-- Copyright (C) 2020  Intel Corporation. All rights reserved.
-- Your use of Intel Corporation's design tools, logic functions 
-- and other software and tools, and any partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Intel Program License 
-- Subscription Agreement, the Intel Quartus Prime License Agreement,
-- the Intel FPGA IP License Agreement, or other applicable license
-- agreement, including, without limitation, that your use is for
-- the sole purpose of programming logic devices manufactured by
-- Intel and sold by Intel or its authorized distributors.  Please
-- refer to the applicable agreement for further details, at
-- https://fpgasoftware.intel.com/eula.

-- PROGRAM		"Quartus Prime"
-- VERSION		"Version 20.1.0 Build 711 06/05/2020 SJ Lite Edition"
-- CREATED		"Thu Nov 12 15:51:03 2020"

LIBRARY ieee;
USE ieee.std_logic_1164.all; 

LIBRARY work;

ENTITY alucontrol IS 
	PORT
	(
		AluOP :  IN  STD_LOGIC_VECTOR(1 DOWNTO 0);
		FunctionInput :  IN  STD_LOGIC_VECTOR(5 DOWNTO 0);
		AluControlFunction :  OUT  STD_LOGIC_VECTOR(3 DOWNTO 0)
	);
END alucontrol;

ARCHITECTURE bdf_type OF alucontrol IS 

SIGNAL	AluControlFunction_ALTERA_SYNTHESIZED :  STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_61 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_62 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_63 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_64 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_65 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_66 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_67 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_68 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_9 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_10 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_17 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_18 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_69 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_25 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_70 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_71 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_72 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_73 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_74 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_75 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_76 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_41 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_77 :  STD_LOGIC;


BEGIN 



SYNTHESIZED_WIRE_62 <= NOT(AluOP(1));



SYNTHESIZED_WIRE_74 <= NOT(SYNTHESIZED_WIRE_61);



SYNTHESIZED_WIRE_10 <= SYNTHESIZED_WIRE_62 AND SYNTHESIZED_WIRE_63;


SYNTHESIZED_WIRE_9 <= AluOP(1) AND FunctionInput(5) AND SYNTHESIZED_WIRE_63 AND SYNTHESIZED_WIRE_64 AND SYNTHESIZED_WIRE_65 AND SYNTHESIZED_WIRE_66 AND SYNTHESIZED_WIRE_67 AND SYNTHESIZED_WIRE_68;


SYNTHESIZED_WIRE_77 <= SYNTHESIZED_WIRE_9 OR SYNTHESIZED_WIRE_10;


SYNTHESIZED_WIRE_18 <= SYNTHESIZED_WIRE_62 AND AluOP(0);


SYNTHESIZED_WIRE_17 <= AluOP(1) AND FunctionInput(5) AND SYNTHESIZED_WIRE_63 AND SYNTHESIZED_WIRE_64 AND FunctionInput(1) AND SYNTHESIZED_WIRE_66 AND SYNTHESIZED_WIRE_67 AND SYNTHESIZED_WIRE_68;


SYNTHESIZED_WIRE_61 <= SYNTHESIZED_WIRE_17 OR SYNTHESIZED_WIRE_18;


SYNTHESIZED_WIRE_69 <= AluOP(1) AND AluOP(0);


SYNTHESIZED_WIRE_73 <= NOT(SYNTHESIZED_WIRE_69);



SYNTHESIZED_WIRE_25 <= AluOP(1) AND FunctionInput(5) AND SYNTHESIZED_WIRE_63 AND SYNTHESIZED_WIRE_64 AND SYNTHESIZED_WIRE_65 AND FunctionInput(2) AND SYNTHESIZED_WIRE_67 AND SYNTHESIZED_WIRE_68;


SYNTHESIZED_WIRE_63 <= NOT(AluOP(0));



SYNTHESIZED_WIRE_75 <= NOT(SYNTHESIZED_WIRE_25);



SYNTHESIZED_WIRE_70 <= AluOP(1) AND FunctionInput(5) AND SYNTHESIZED_WIRE_63 AND SYNTHESIZED_WIRE_64 AND SYNTHESIZED_WIRE_65 AND FunctionInput(2) AND FunctionInput(0) AND SYNTHESIZED_WIRE_68;


SYNTHESIZED_WIRE_76 <= NOT(SYNTHESIZED_WIRE_70);



SYNTHESIZED_WIRE_71 <= AluOP(1) AND FunctionInput(5) AND SYNTHESIZED_WIRE_63 AND SYNTHESIZED_WIRE_64 AND FunctionInput(1) AND SYNTHESIZED_WIRE_66 AND SYNTHESIZED_WIRE_67 AND FunctionInput(3);


SYNTHESIZED_WIRE_41 <= NOT(SYNTHESIZED_WIRE_71);



AluControlFunction_ALTERA_SYNTHESIZED(3) <= SYNTHESIZED_WIRE_72 OR SYNTHESIZED_WIRE_73 OR SYNTHESIZED_WIRE_74 OR SYNTHESIZED_WIRE_75 OR SYNTHESIZED_WIRE_76 OR SYNTHESIZED_WIRE_41;


AluControlFunction_ALTERA_SYNTHESIZED(2) <= SYNTHESIZED_WIRE_72 OR SYNTHESIZED_WIRE_75 OR SYNTHESIZED_WIRE_73 OR SYNTHESIZED_WIRE_76 OR SYNTHESIZED_WIRE_71 OR SYNTHESIZED_WIRE_61;


AluControlFunction_ALTERA_SYNTHESIZED(1) <= SYNTHESIZED_WIRE_77 OR SYNTHESIZED_WIRE_69 OR SYNTHESIZED_WIRE_61 OR SYNTHESIZED_WIRE_75 OR SYNTHESIZED_WIRE_76 OR SYNTHESIZED_WIRE_71;


AluControlFunction_ALTERA_SYNTHESIZED(0) <= SYNTHESIZED_WIRE_72 OR SYNTHESIZED_WIRE_69 OR SYNTHESIZED_WIRE_74 OR SYNTHESIZED_WIRE_75 OR SYNTHESIZED_WIRE_70 OR SYNTHESIZED_WIRE_71;



SYNTHESIZED_WIRE_64 <= NOT(FunctionInput(4));



SYNTHESIZED_WIRE_68 <= NOT(FunctionInput(3));



SYNTHESIZED_WIRE_66 <= NOT(FunctionInput(2));



SYNTHESIZED_WIRE_65 <= NOT(FunctionInput(1));



SYNTHESIZED_WIRE_67 <= NOT(FunctionInput(0));



SYNTHESIZED_WIRE_72 <= NOT(SYNTHESIZED_WIRE_77);


AluControlFunction <= AluControlFunction_ALTERA_SYNTHESIZED;

END bdf_type;