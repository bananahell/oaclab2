-- Copyright (C) 2020  Intel Corporation. All rights reserved.
-- Your use of Intel Corporation's design tools, logic functions 
-- and other software and tools, and any partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Intel Program License 
-- Subscription Agreement, the Intel Quartus Prime License Agreement,
-- the Intel FPGA IP License Agreement, or other applicable license
-- agreement, including, without limitation, that your use is for
-- the sole purpose of programming logic devices manufactured by
-- Intel and sold by Intel or its authorized distributors.  Please
-- refer to the applicable agreement for further details, at
-- https://fpgasoftware.intel.com/eula.

-- PROGRAM		"Quartus Prime"
-- VERSION		"Version 20.1.0 Build 711 06/05/2020 SJ Lite Edition"
-- CREATED		"Thu Nov 12 18:01:21 2020"

LIBRARY ieee;
USE ieee.std_logic_1164.all; 

LIBRARY work;

ENTITY \32writeenabledflipflop32bit\ IS 
	PORT
	(
		WriteEnable :  IN  STD_LOGIC;
		ClockInput :  IN  STD_LOGIC;
		Input :  IN  STD_LOGIC_VECTOR(31 DOWNTO 0);
		Selector :  IN  STD_LOGIC_VECTOR(0 TO 4);
		ResultPin :  OUT  STD_LOGIC_VECTOR(31 DOWNTO 0)
	);
END \32writeenabledflipflop32bit\;

ARCHITECTURE bdf_type OF \32writeenabledflipflop32bit\ IS 

COMPONENT mux32_32bit
	PORT(Input00 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 Input01 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 Input02 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 Input03 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 Input04 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 Input05 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 Input06 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 Input07 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 Input08 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 Input09 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 Input10 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 Input11 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 Input12 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 Input13 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 Input14 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 Input15 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 Input16 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 Input17 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 Input18 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 Input19 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 Input20 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 Input21 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 Input22 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 Input23 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 Input24 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 Input25 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 Input26 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 Input27 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 Input28 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 Input29 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 Input30 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 Input31 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 Selector : IN STD_LOGIC_VECTOR(4 DOWNTO 0);
		 ResultPin : OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
	);
END COMPONENT;

COMPONENT writeenabledflipflop32bit
	PORT(WriteEnable : IN STD_LOGIC;
		 ClockInput : IN STD_LOGIC;
		 Input : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 OutputRes : OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
	);
END COMPONENT;

COMPONENT and5_1bit
	PORT(Input1 : IN STD_LOGIC;
		 Input2 : IN STD_LOGIC;
		 Input3 : IN STD_LOGIC;
		 Input5 : IN STD_LOGIC;
		 Input4 : IN STD_LOGIC;
		 ResultingPin : OUT STD_LOGIC
	);
END COMPONENT;

SIGNAL	SYNTHESIZED_WIRE_0 :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_1 :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_2 :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_3 :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_4 :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_5 :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_6 :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_7 :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_8 :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_9 :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_10 :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_11 :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_12 :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_13 :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_14 :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_15 :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_16 :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_17 :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_18 :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_19 :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_20 :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_21 :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_22 :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_23 :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_24 :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_25 :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_26 :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_27 :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_28 :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_29 :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_30 :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_31 :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_32 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_33 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_34 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_35 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_36 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_37 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_38 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_39 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_40 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_41 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_42 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_43 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_44 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_45 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_46 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_47 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_48 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_49 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_50 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_51 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_52 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_53 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_54 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_55 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_56 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_57 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_58 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_59 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_60 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_61 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_62 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_63 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_64 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_65 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_66 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_67 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_68 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_69 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_70 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_71 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_72 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_73 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_74 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_75 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_76 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_77 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_78 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_79 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_80 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_81 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_82 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_83 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_84 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_85 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_86 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_87 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_88 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_89 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_90 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_91 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_92 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_93 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_94 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_95 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_96 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_97 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_98 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_99 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_100 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_101 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_102 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_103 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_104 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_105 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_106 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_107 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_108 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_109 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_110 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_111 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_112 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_113 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_114 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_115 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_116 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_117 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_118 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_119 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_120 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_121 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_122 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_123 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_124 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_125 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_126 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_127 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_128 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_129 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_130 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_131 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_132 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_133 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_134 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_135 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_136 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_137 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_138 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_139 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_140 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_141 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_142 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_143 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_144 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_145 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_146 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_147 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_148 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_149 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_150 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_151 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_152 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_153 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_154 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_155 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_156 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_157 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_158 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_159 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_160 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_161 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_162 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_163 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_164 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_165 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_166 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_167 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_168 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_169 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_170 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_171 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_172 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_173 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_174 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_175 :  STD_LOGIC;


BEGIN 



b2v_inst : mux32_32bit
PORT MAP(Input00 => SYNTHESIZED_WIRE_0,
		 Input01 => SYNTHESIZED_WIRE_1,
		 Input02 => SYNTHESIZED_WIRE_2,
		 Input03 => SYNTHESIZED_WIRE_3,
		 Input04 => SYNTHESIZED_WIRE_4,
		 Input05 => SYNTHESIZED_WIRE_5,
		 Input06 => SYNTHESIZED_WIRE_6,
		 Input07 => SYNTHESIZED_WIRE_7,
		 Input08 => SYNTHESIZED_WIRE_8,
		 Input09 => SYNTHESIZED_WIRE_9,
		 Input10 => SYNTHESIZED_WIRE_10,
		 Input11 => SYNTHESIZED_WIRE_11,
		 Input12 => SYNTHESIZED_WIRE_12,
		 Input13 => SYNTHESIZED_WIRE_13,
		 Input14 => SYNTHESIZED_WIRE_14,
		 Input15 => SYNTHESIZED_WIRE_15,
		 Input16 => SYNTHESIZED_WIRE_16,
		 Input17 => SYNTHESIZED_WIRE_17,
		 Input18 => SYNTHESIZED_WIRE_18,
		 Input19 => SYNTHESIZED_WIRE_19,
		 Input20 => SYNTHESIZED_WIRE_20,
		 Input21 => SYNTHESIZED_WIRE_21,
		 Input22 => SYNTHESIZED_WIRE_22,
		 Input23 => SYNTHESIZED_WIRE_23,
		 Input24 => SYNTHESIZED_WIRE_24,
		 Input25 => SYNTHESIZED_WIRE_25,
		 Input26 => SYNTHESIZED_WIRE_26,
		 Input27 => SYNTHESIZED_WIRE_27,
		 Input28 => SYNTHESIZED_WIRE_28,
		 Input29 => SYNTHESIZED_WIRE_29,
		 Input30 => SYNTHESIZED_WIRE_30,
		 Input31 => SYNTHESIZED_WIRE_31,
		 Selector => Selector,
		 ResultPin => ResultPin);


SYNTHESIZED_WIRE_104 <= NOT(Selector(4));



SYNTHESIZED_WIRE_100 <= NOT(Selector(4));



SYNTHESIZED_WIRE_101 <= NOT(Selector(3));



SYNTHESIZED_WIRE_64 <= SYNTHESIZED_WIRE_32 AND ClockInput;


SYNTHESIZED_WIRE_65 <= SYNTHESIZED_WIRE_33 AND ClockInput;


SYNTHESIZED_WIRE_66 <= SYNTHESIZED_WIRE_34 AND ClockInput;


SYNTHESIZED_WIRE_67 <= SYNTHESIZED_WIRE_35 AND ClockInput;


SYNTHESIZED_WIRE_68 <= SYNTHESIZED_WIRE_36 AND ClockInput;


SYNTHESIZED_WIRE_69 <= SYNTHESIZED_WIRE_37 AND ClockInput;


SYNTHESIZED_WIRE_70 <= SYNTHESIZED_WIRE_38 AND ClockInput;


SYNTHESIZED_WIRE_102 <= NOT(Selector(2));



SYNTHESIZED_WIRE_71 <= SYNTHESIZED_WIRE_39 AND ClockInput;


SYNTHESIZED_WIRE_72 <= SYNTHESIZED_WIRE_40 AND ClockInput;


SYNTHESIZED_WIRE_73 <= SYNTHESIZED_WIRE_41 AND ClockInput;


SYNTHESIZED_WIRE_74 <= SYNTHESIZED_WIRE_42 AND ClockInput;


SYNTHESIZED_WIRE_75 <= SYNTHESIZED_WIRE_43 AND ClockInput;


SYNTHESIZED_WIRE_76 <= SYNTHESIZED_WIRE_44 AND ClockInput;


SYNTHESIZED_WIRE_77 <= SYNTHESIZED_WIRE_45 AND ClockInput;


SYNTHESIZED_WIRE_78 <= SYNTHESIZED_WIRE_46 AND ClockInput;


SYNTHESIZED_WIRE_79 <= SYNTHESIZED_WIRE_47 AND ClockInput;


SYNTHESIZED_WIRE_80 <= SYNTHESIZED_WIRE_48 AND ClockInput;


SYNTHESIZED_WIRE_103 <= NOT(Selector(0));



SYNTHESIZED_WIRE_81 <= SYNTHESIZED_WIRE_49 AND ClockInput;


SYNTHESIZED_WIRE_82 <= SYNTHESIZED_WIRE_50 AND ClockInput;


SYNTHESIZED_WIRE_83 <= SYNTHESIZED_WIRE_51 AND ClockInput;


SYNTHESIZED_WIRE_84 <= SYNTHESIZED_WIRE_52 AND ClockInput;


SYNTHESIZED_WIRE_85 <= SYNTHESIZED_WIRE_53 AND ClockInput;


SYNTHESIZED_WIRE_86 <= SYNTHESIZED_WIRE_54 AND ClockInput;


SYNTHESIZED_WIRE_87 <= SYNTHESIZED_WIRE_55 AND ClockInput;


SYNTHESIZED_WIRE_88 <= SYNTHESIZED_WIRE_56 AND ClockInput;


SYNTHESIZED_WIRE_89 <= SYNTHESIZED_WIRE_57 AND ClockInput;


SYNTHESIZED_WIRE_90 <= SYNTHESIZED_WIRE_58 AND ClockInput;


SYNTHESIZED_WIRE_109 <= NOT(Selector(4));



SYNTHESIZED_WIRE_91 <= SYNTHESIZED_WIRE_59 AND ClockInput;


SYNTHESIZED_WIRE_92 <= SYNTHESIZED_WIRE_60 AND ClockInput;


SYNTHESIZED_WIRE_93 <= SYNTHESIZED_WIRE_61 AND ClockInput;


SYNTHESIZED_WIRE_94 <= SYNTHESIZED_WIRE_62 AND ClockInput;


SYNTHESIZED_WIRE_95 <= SYNTHESIZED_WIRE_63 AND ClockInput;


b2v_inst145 : writeenabledflipflop32bit
PORT MAP(WriteEnable => WriteEnable,
		 ClockInput => SYNTHESIZED_WIRE_64,
		 Input => Input,
		 OutputRes => SYNTHESIZED_WIRE_0);


b2v_inst146 : writeenabledflipflop32bit
PORT MAP(WriteEnable => WriteEnable,
		 ClockInput => SYNTHESIZED_WIRE_65,
		 Input => Input,
		 OutputRes => SYNTHESIZED_WIRE_1);


b2v_inst147 : writeenabledflipflop32bit
PORT MAP(WriteEnable => WriteEnable,
		 ClockInput => SYNTHESIZED_WIRE_66,
		 Input => Input,
		 OutputRes => SYNTHESIZED_WIRE_2);


b2v_inst148 : writeenabledflipflop32bit
PORT MAP(WriteEnable => WriteEnable,
		 ClockInput => SYNTHESIZED_WIRE_67,
		 Input => Input,
		 OutputRes => SYNTHESIZED_WIRE_3);


b2v_inst149 : writeenabledflipflop32bit
PORT MAP(WriteEnable => WriteEnable,
		 ClockInput => SYNTHESIZED_WIRE_68,
		 Input => Input,
		 OutputRes => SYNTHESIZED_WIRE_4);


SYNTHESIZED_WIRE_110 <= NOT(Selector(3));



b2v_inst150 : writeenabledflipflop32bit
PORT MAP(WriteEnable => WriteEnable,
		 ClockInput => SYNTHESIZED_WIRE_69,
		 Input => Input,
		 OutputRes => SYNTHESIZED_WIRE_5);


b2v_inst151 : writeenabledflipflop32bit
PORT MAP(WriteEnable => WriteEnable,
		 ClockInput => SYNTHESIZED_WIRE_70,
		 Input => Input,
		 OutputRes => SYNTHESIZED_WIRE_6);


b2v_inst152 : writeenabledflipflop32bit
PORT MAP(WriteEnable => WriteEnable,
		 ClockInput => SYNTHESIZED_WIRE_71,
		 Input => Input,
		 OutputRes => SYNTHESIZED_WIRE_7);


b2v_inst153 : writeenabledflipflop32bit
PORT MAP(WriteEnable => WriteEnable,
		 ClockInput => SYNTHESIZED_WIRE_72,
		 Input => Input,
		 OutputRes => SYNTHESIZED_WIRE_8);


b2v_inst154 : writeenabledflipflop32bit
PORT MAP(WriteEnable => WriteEnable,
		 ClockInput => SYNTHESIZED_WIRE_73,
		 Input => Input,
		 OutputRes => SYNTHESIZED_WIRE_9);


b2v_inst155 : writeenabledflipflop32bit
PORT MAP(WriteEnable => WriteEnable,
		 ClockInput => SYNTHESIZED_WIRE_74,
		 Input => Input,
		 OutputRes => SYNTHESIZED_WIRE_10);


b2v_inst156 : writeenabledflipflop32bit
PORT MAP(WriteEnable => WriteEnable,
		 ClockInput => SYNTHESIZED_WIRE_75,
		 Input => Input,
		 OutputRes => SYNTHESIZED_WIRE_11);


b2v_inst157 : writeenabledflipflop32bit
PORT MAP(WriteEnable => WriteEnable,
		 ClockInput => SYNTHESIZED_WIRE_76,
		 Input => Input,
		 OutputRes => SYNTHESIZED_WIRE_12);


b2v_inst158 : writeenabledflipflop32bit
PORT MAP(WriteEnable => WriteEnable,
		 ClockInput => SYNTHESIZED_WIRE_77,
		 Input => Input,
		 OutputRes => SYNTHESIZED_WIRE_13);


b2v_inst159 : writeenabledflipflop32bit
PORT MAP(WriteEnable => WriteEnable,
		 ClockInput => SYNTHESIZED_WIRE_78,
		 Input => Input,
		 OutputRes => SYNTHESIZED_WIRE_14);


SYNTHESIZED_WIRE_111 <= NOT(Selector(2));



b2v_inst160 : writeenabledflipflop32bit
PORT MAP(WriteEnable => WriteEnable,
		 ClockInput => SYNTHESIZED_WIRE_79,
		 Input => Input,
		 OutputRes => SYNTHESIZED_WIRE_15);


b2v_inst161 : writeenabledflipflop32bit
PORT MAP(WriteEnable => WriteEnable,
		 ClockInput => SYNTHESIZED_WIRE_80,
		 Input => Input,
		 OutputRes => SYNTHESIZED_WIRE_16);


b2v_inst162 : writeenabledflipflop32bit
PORT MAP(WriteEnable => WriteEnable,
		 ClockInput => SYNTHESIZED_WIRE_81,
		 Input => Input,
		 OutputRes => SYNTHESIZED_WIRE_17);


b2v_inst163 : writeenabledflipflop32bit
PORT MAP(WriteEnable => WriteEnable,
		 ClockInput => SYNTHESIZED_WIRE_82,
		 Input => Input,
		 OutputRes => SYNTHESIZED_WIRE_18);


b2v_inst164 : writeenabledflipflop32bit
PORT MAP(WriteEnable => WriteEnable,
		 ClockInput => SYNTHESIZED_WIRE_83,
		 Input => Input,
		 OutputRes => SYNTHESIZED_WIRE_19);


b2v_inst165 : writeenabledflipflop32bit
PORT MAP(WriteEnable => WriteEnable,
		 ClockInput => SYNTHESIZED_WIRE_84,
		 Input => Input,
		 OutputRes => SYNTHESIZED_WIRE_20);


b2v_inst166 : writeenabledflipflop32bit
PORT MAP(WriteEnable => WriteEnable,
		 ClockInput => SYNTHESIZED_WIRE_85,
		 Input => Input,
		 OutputRes => SYNTHESIZED_WIRE_21);


b2v_inst167 : writeenabledflipflop32bit
PORT MAP(WriteEnable => WriteEnable,
		 ClockInput => SYNTHESIZED_WIRE_86,
		 Input => Input,
		 OutputRes => SYNTHESIZED_WIRE_22);


b2v_inst168 : writeenabledflipflop32bit
PORT MAP(WriteEnable => WriteEnable,
		 ClockInput => SYNTHESIZED_WIRE_87,
		 Input => Input,
		 OutputRes => SYNTHESIZED_WIRE_23);


b2v_inst169 : writeenabledflipflop32bit
PORT MAP(WriteEnable => WriteEnable,
		 ClockInput => SYNTHESIZED_WIRE_88,
		 Input => Input,
		 OutputRes => SYNTHESIZED_WIRE_24);


SYNTHESIZED_WIRE_117 <= NOT(Selector(4));



b2v_inst170 : writeenabledflipflop32bit
PORT MAP(WriteEnable => WriteEnable,
		 ClockInput => SYNTHESIZED_WIRE_89,
		 Input => Input,
		 OutputRes => SYNTHESIZED_WIRE_25);


b2v_inst171 : writeenabledflipflop32bit
PORT MAP(WriteEnable => WriteEnable,
		 ClockInput => SYNTHESIZED_WIRE_90,
		 Input => Input,
		 OutputRes => SYNTHESIZED_WIRE_26);


b2v_inst172 : writeenabledflipflop32bit
PORT MAP(WriteEnable => WriteEnable,
		 ClockInput => SYNTHESIZED_WIRE_91,
		 Input => Input,
		 OutputRes => SYNTHESIZED_WIRE_27);


b2v_inst173 : writeenabledflipflop32bit
PORT MAP(WriteEnable => WriteEnable,
		 ClockInput => SYNTHESIZED_WIRE_92,
		 Input => Input,
		 OutputRes => SYNTHESIZED_WIRE_28);


b2v_inst174 : writeenabledflipflop32bit
PORT MAP(WriteEnable => WriteEnable,
		 ClockInput => SYNTHESIZED_WIRE_93,
		 Input => Input,
		 OutputRes => SYNTHESIZED_WIRE_29);


b2v_inst175 : writeenabledflipflop32bit
PORT MAP(WriteEnable => WriteEnable,
		 ClockInput => SYNTHESIZED_WIRE_94,
		 Input => Input,
		 OutputRes => SYNTHESIZED_WIRE_30);


b2v_inst176 : writeenabledflipflop32bit
PORT MAP(WriteEnable => WriteEnable,
		 ClockInput => SYNTHESIZED_WIRE_95,
		 Input => Input,
		 OutputRes => SYNTHESIZED_WIRE_31);


SYNTHESIZED_WIRE_118 <= NOT(Selector(3));



b2v_inst183 : and5_1bit
PORT MAP(Input1 => SYNTHESIZED_WIRE_96,
		 Input2 => SYNTHESIZED_WIRE_97,
		 Input3 => SYNTHESIZED_WIRE_98,
		 Input5 => SYNTHESIZED_WIRE_99,
		 Input4 => Selector(0),
		 ResultingPin => SYNTHESIZED_WIRE_33);


b2v_inst184 : and5_1bit
PORT MAP(Input1 => SYNTHESIZED_WIRE_100,
		 Input2 => SYNTHESIZED_WIRE_101,
		 Input3 => SYNTHESIZED_WIRE_102,
		 Input5 => Selector(1),
		 Input4 => SYNTHESIZED_WIRE_103,
		 ResultingPin => SYNTHESIZED_WIRE_34);


b2v_inst185 : and5_1bit
PORT MAP(Input1 => SYNTHESIZED_WIRE_104,
		 Input2 => SYNTHESIZED_WIRE_105,
		 Input3 => SYNTHESIZED_WIRE_106,
		 Input5 => SYNTHESIZED_WIRE_107,
		 Input4 => SYNTHESIZED_WIRE_108,
		 ResultingPin => SYNTHESIZED_WIRE_32);


b2v_inst186 : and5_1bit
PORT MAP(Input1 => SYNTHESIZED_WIRE_109,
		 Input2 => SYNTHESIZED_WIRE_110,
		 Input3 => SYNTHESIZED_WIRE_111,
		 Input5 => Selector(1),
		 Input4 => Selector(0),
		 ResultingPin => SYNTHESIZED_WIRE_35);


b2v_inst187 : and5_1bit
PORT MAP(Input1 => SYNTHESIZED_WIRE_112,
		 Input2 => SYNTHESIZED_WIRE_113,
		 Input3 => Selector(2),
		 Input5 => Selector(1),
		 Input4 => SYNTHESIZED_WIRE_114,
		 ResultingPin => SYNTHESIZED_WIRE_38);


b2v_inst188 : and5_1bit
PORT MAP(Input1 => SYNTHESIZED_WIRE_115,
		 Input2 => SYNTHESIZED_WIRE_116,
		 Input3 => Selector(2),
		 Input5 => Selector(1),
		 Input4 => Selector(0),
		 ResultingPin => SYNTHESIZED_WIRE_39);


b2v_inst189 : and5_1bit
PORT MAP(Input1 => SYNTHESIZED_WIRE_117,
		 Input2 => SYNTHESIZED_WIRE_118,
		 Input3 => Selector(2),
		 Input5 => SYNTHESIZED_WIRE_119,
		 Input4 => SYNTHESIZED_WIRE_120,
		 ResultingPin => SYNTHESIZED_WIRE_36);


SYNTHESIZED_WIRE_119 <= NOT(Selector(1));



b2v_inst190 : and5_1bit
PORT MAP(Input1 => SYNTHESIZED_WIRE_121,
		 Input2 => SYNTHESIZED_WIRE_122,
		 Input3 => Selector(2),
		 Input5 => SYNTHESIZED_WIRE_123,
		 Input4 => Selector(0),
		 ResultingPin => SYNTHESIZED_WIRE_37);


b2v_inst191 : and5_1bit
PORT MAP(Input1 => SYNTHESIZED_WIRE_124,
		 Input2 => Selector(3),
		 Input3 => SYNTHESIZED_WIRE_125,
		 Input5 => SYNTHESIZED_WIRE_126,
		 Input4 => SYNTHESIZED_WIRE_127,
		 ResultingPin => SYNTHESIZED_WIRE_40);


b2v_inst192 : and5_1bit
PORT MAP(Input1 => SYNTHESIZED_WIRE_128,
		 Input2 => Selector(3),
		 Input3 => SYNTHESIZED_WIRE_129,
		 Input5 => SYNTHESIZED_WIRE_130,
		 Input4 => Selector(0),
		 ResultingPin => SYNTHESIZED_WIRE_41);


b2v_inst193 : and5_1bit
PORT MAP(Input1 => SYNTHESIZED_WIRE_131,
		 Input2 => Selector(3),
		 Input3 => SYNTHESIZED_WIRE_132,
		 Input5 => Selector(1),
		 Input4 => SYNTHESIZED_WIRE_133,
		 ResultingPin => SYNTHESIZED_WIRE_42);


b2v_inst194 : and5_1bit
PORT MAP(Input1 => SYNTHESIZED_WIRE_134,
		 Input2 => Selector(3),
		 Input3 => SYNTHESIZED_WIRE_135,
		 Input5 => Selector(1),
		 Input4 => Selector(0),
		 ResultingPin => SYNTHESIZED_WIRE_43);


b2v_inst195 : and5_1bit
PORT MAP(Input1 => SYNTHESIZED_WIRE_136,
		 Input2 => Selector(3),
		 Input3 => Selector(2),
		 Input5 => SYNTHESIZED_WIRE_137,
		 Input4 => SYNTHESIZED_WIRE_138,
		 ResultingPin => SYNTHESIZED_WIRE_44);


b2v_inst196 : and5_1bit
PORT MAP(Input1 => SYNTHESIZED_WIRE_139,
		 Input2 => Selector(3),
		 Input3 => Selector(2),
		 Input5 => SYNTHESIZED_WIRE_140,
		 Input4 => Selector(0),
		 ResultingPin => SYNTHESIZED_WIRE_45);


b2v_inst197 : and5_1bit
PORT MAP(Input1 => SYNTHESIZED_WIRE_141,
		 Input2 => Selector(3),
		 Input3 => Selector(2),
		 Input5 => Selector(1),
		 Input4 => SYNTHESIZED_WIRE_142,
		 ResultingPin => SYNTHESIZED_WIRE_46);


b2v_inst198 : and5_1bit
PORT MAP(Input1 => SYNTHESIZED_WIRE_143,
		 Input2 => Selector(3),
		 Input3 => Selector(2),
		 Input5 => Selector(1),
		 Input4 => Selector(0),
		 ResultingPin => SYNTHESIZED_WIRE_47);


b2v_inst199 : and5_1bit
PORT MAP(Input1 => Selector(4),
		 Input2 => SYNTHESIZED_WIRE_144,
		 Input3 => SYNTHESIZED_WIRE_145,
		 Input5 => SYNTHESIZED_WIRE_146,
		 Input4 => SYNTHESIZED_WIRE_147,
		 ResultingPin => SYNTHESIZED_WIRE_48);


SYNTHESIZED_WIRE_105 <= NOT(Selector(3));



SYNTHESIZED_WIRE_120 <= NOT(Selector(0));



b2v_inst200 : and5_1bit
PORT MAP(Input1 => Selector(4),
		 Input2 => SYNTHESIZED_WIRE_148,
		 Input3 => SYNTHESIZED_WIRE_149,
		 Input5 => SYNTHESIZED_WIRE_150,
		 Input4 => Selector(0),
		 ResultingPin => SYNTHESIZED_WIRE_49);


b2v_inst201 : and5_1bit
PORT MAP(Input1 => Selector(4),
		 Input2 => SYNTHESIZED_WIRE_151,
		 Input3 => SYNTHESIZED_WIRE_152,
		 Input5 => Selector(1),
		 Input4 => SYNTHESIZED_WIRE_153,
		 ResultingPin => SYNTHESIZED_WIRE_50);


b2v_inst202 : and5_1bit
PORT MAP(Input1 => Selector(4),
		 Input2 => SYNTHESIZED_WIRE_154,
		 Input3 => SYNTHESIZED_WIRE_155,
		 Input5 => Selector(1),
		 Input4 => Selector(0),
		 ResultingPin => SYNTHESIZED_WIRE_51);


b2v_inst203 : and5_1bit
PORT MAP(Input1 => Selector(4),
		 Input2 => SYNTHESIZED_WIRE_156,
		 Input3 => Selector(2),
		 Input5 => SYNTHESIZED_WIRE_157,
		 Input4 => SYNTHESIZED_WIRE_158,
		 ResultingPin => SYNTHESIZED_WIRE_52);


b2v_inst204 : and5_1bit
PORT MAP(Input1 => Selector(4),
		 Input2 => SYNTHESIZED_WIRE_159,
		 Input3 => Selector(2),
		 Input5 => SYNTHESIZED_WIRE_160,
		 Input4 => Selector(0),
		 ResultingPin => SYNTHESIZED_WIRE_53);


b2v_inst205 : and5_1bit
PORT MAP(Input1 => Selector(4),
		 Input2 => SYNTHESIZED_WIRE_161,
		 Input3 => Selector(2),
		 Input5 => Selector(1),
		 Input4 => SYNTHESIZED_WIRE_162,
		 ResultingPin => SYNTHESIZED_WIRE_54);


b2v_inst206 : and5_1bit
PORT MAP(Input1 => Selector(4),
		 Input2 => SYNTHESIZED_WIRE_163,
		 Input3 => Selector(2),
		 Input5 => Selector(1),
		 Input4 => Selector(0),
		 ResultingPin => SYNTHESIZED_WIRE_55);


b2v_inst207 : and5_1bit
PORT MAP(Input1 => Selector(4),
		 Input2 => Selector(3),
		 Input3 => SYNTHESIZED_WIRE_164,
		 Input5 => SYNTHESIZED_WIRE_165,
		 Input4 => SYNTHESIZED_WIRE_166,
		 ResultingPin => SYNTHESIZED_WIRE_56);


b2v_inst208 : and5_1bit
PORT MAP(Input1 => Selector(4),
		 Input2 => Selector(3),
		 Input3 => SYNTHESIZED_WIRE_167,
		 Input5 => SYNTHESIZED_WIRE_168,
		 Input4 => Selector(0),
		 ResultingPin => SYNTHESIZED_WIRE_57);


b2v_inst209 : and5_1bit
PORT MAP(Input1 => Selector(4),
		 Input2 => Selector(3),
		 Input3 => SYNTHESIZED_WIRE_169,
		 Input5 => Selector(1),
		 Input4 => SYNTHESIZED_WIRE_170,
		 ResultingPin => SYNTHESIZED_WIRE_58);


SYNTHESIZED_WIRE_121 <= NOT(Selector(4));



b2v_inst210 : and5_1bit
PORT MAP(Input1 => Selector(4),
		 Input2 => Selector(3),
		 Input3 => SYNTHESIZED_WIRE_171,
		 Input5 => Selector(1),
		 Input4 => Selector(0),
		 ResultingPin => SYNTHESIZED_WIRE_59);


b2v_inst211 : and5_1bit
PORT MAP(Input1 => Selector(4),
		 Input2 => Selector(3),
		 Input3 => Selector(2),
		 Input5 => SYNTHESIZED_WIRE_172,
		 Input4 => SYNTHESIZED_WIRE_173,
		 ResultingPin => SYNTHESIZED_WIRE_60);


b2v_inst212 : and5_1bit
PORT MAP(Input1 => Selector(4),
		 Input2 => Selector(3),
		 Input3 => Selector(2),
		 Input5 => SYNTHESIZED_WIRE_174,
		 Input4 => Selector(0),
		 ResultingPin => SYNTHESIZED_WIRE_61);


b2v_inst213 : and5_1bit
PORT MAP(Input1 => Selector(4),
		 Input2 => Selector(3),
		 Input3 => Selector(2),
		 Input5 => Selector(1),
		 Input4 => SYNTHESIZED_WIRE_175,
		 ResultingPin => SYNTHESIZED_WIRE_62);


b2v_inst214 : and5_1bit
PORT MAP(Input1 => Selector(4),
		 Input2 => Selector(3),
		 Input3 => Selector(2),
		 Input5 => Selector(1),
		 Input4 => Selector(0),
		 ResultingPin => SYNTHESIZED_WIRE_63);


SYNTHESIZED_WIRE_122 <= NOT(Selector(3));



SYNTHESIZED_WIRE_123 <= NOT(Selector(1));



SYNTHESIZED_WIRE_112 <= NOT(Selector(4));



SYNTHESIZED_WIRE_113 <= NOT(Selector(3));



SYNTHESIZED_WIRE_114 <= NOT(Selector(0));



SYNTHESIZED_WIRE_115 <= NOT(Selector(4));



SYNTHESIZED_WIRE_116 <= NOT(Selector(3));



SYNTHESIZED_WIRE_124 <= NOT(Selector(4));



SYNTHESIZED_WIRE_106 <= NOT(Selector(2));



SYNTHESIZED_WIRE_125 <= NOT(Selector(2));



SYNTHESIZED_WIRE_126 <= NOT(Selector(1));



SYNTHESIZED_WIRE_127 <= NOT(Selector(0));



SYNTHESIZED_WIRE_128 <= NOT(Selector(4));



SYNTHESIZED_WIRE_129 <= NOT(Selector(2));



SYNTHESIZED_WIRE_130 <= NOT(Selector(1));



SYNTHESIZED_WIRE_131 <= NOT(Selector(4));



SYNTHESIZED_WIRE_132 <= NOT(Selector(2));



SYNTHESIZED_WIRE_133 <= NOT(Selector(0));



SYNTHESIZED_WIRE_134 <= NOT(Selector(4));



SYNTHESIZED_WIRE_107 <= NOT(Selector(1));



SYNTHESIZED_WIRE_135 <= NOT(Selector(2));



SYNTHESIZED_WIRE_136 <= NOT(Selector(4));



SYNTHESIZED_WIRE_137 <= NOT(Selector(1));



SYNTHESIZED_WIRE_138 <= NOT(Selector(0));



SYNTHESIZED_WIRE_139 <= NOT(Selector(4));



SYNTHESIZED_WIRE_140 <= NOT(Selector(1));



SYNTHESIZED_WIRE_141 <= NOT(Selector(4));



SYNTHESIZED_WIRE_142 <= NOT(Selector(0));



SYNTHESIZED_WIRE_143 <= NOT(Selector(4));



SYNTHESIZED_WIRE_144 <= NOT(Selector(3));



SYNTHESIZED_WIRE_108 <= NOT(Selector(0));



SYNTHESIZED_WIRE_145 <= NOT(Selector(2));



SYNTHESIZED_WIRE_146 <= NOT(Selector(1));



SYNTHESIZED_WIRE_147 <= NOT(Selector(0));



SYNTHESIZED_WIRE_148 <= NOT(Selector(3));



SYNTHESIZED_WIRE_149 <= NOT(Selector(2));



SYNTHESIZED_WIRE_150 <= NOT(Selector(1));



SYNTHESIZED_WIRE_151 <= NOT(Selector(3));



SYNTHESIZED_WIRE_152 <= NOT(Selector(2));



SYNTHESIZED_WIRE_153 <= NOT(Selector(0));



SYNTHESIZED_WIRE_154 <= NOT(Selector(3));



SYNTHESIZED_WIRE_96 <= NOT(Selector(4));



SYNTHESIZED_WIRE_155 <= NOT(Selector(2));



SYNTHESIZED_WIRE_156 <= NOT(Selector(3));



SYNTHESIZED_WIRE_157 <= NOT(Selector(1));



SYNTHESIZED_WIRE_158 <= NOT(Selector(0));



SYNTHESIZED_WIRE_159 <= NOT(Selector(3));



SYNTHESIZED_WIRE_160 <= NOT(Selector(1));



SYNTHESIZED_WIRE_161 <= NOT(Selector(3));



SYNTHESIZED_WIRE_162 <= NOT(Selector(0));



SYNTHESIZED_WIRE_163 <= NOT(Selector(3));



SYNTHESIZED_WIRE_164 <= NOT(Selector(2));



SYNTHESIZED_WIRE_97 <= NOT(Selector(3));



SYNTHESIZED_WIRE_165 <= NOT(Selector(1));



SYNTHESIZED_WIRE_166 <= NOT(Selector(0));



SYNTHESIZED_WIRE_167 <= NOT(Selector(2));



SYNTHESIZED_WIRE_168 <= NOT(Selector(1));



SYNTHESIZED_WIRE_169 <= NOT(Selector(2));



SYNTHESIZED_WIRE_170 <= NOT(Selector(0));



SYNTHESIZED_WIRE_171 <= NOT(Selector(2));



SYNTHESIZED_WIRE_172 <= NOT(Selector(1));



SYNTHESIZED_WIRE_173 <= NOT(Selector(0));



SYNTHESIZED_WIRE_174 <= NOT(Selector(1));



SYNTHESIZED_WIRE_98 <= NOT(Selector(2));



SYNTHESIZED_WIRE_175 <= NOT(Selector(0));



SYNTHESIZED_WIRE_99 <= NOT(Selector(1));



END bdf_type;