-- Copyright (C) 2020  Intel Corporation. All rights reserved.
-- Your use of Intel Corporation's design tools, logic functions
-- and other software and tools, and any partner logic
-- functions, and any output files from any of the foregoing
-- (including device programming or simulation files), and any
-- associated documentation or information are expressly subject
-- to the terms and conditions of the Intel Program License
-- Subscription Agreement, the Intel Quartus Prime License Agreement,
-- the Intel FPGA IP License Agreement, or other applicable license
-- agreement, including, without limitation, that your use is for
-- the sole purpose of programming logic devices manufactured by
-- Intel and sold by Intel or its authorized distributors.  Please
-- refer to the applicable agreement for further details, at
-- https://fpgasoftware.intel.com/eula.

-- PROGRAM		"Quartus Prime"
-- VERSION		"Version 20.1.0 Build 711 06/05/2020 SJ Lite Edition"
-- CREATED		"Thu Nov 12 18:39:41 2020"

LIBRARY ieee;
USE ieee.std_logic_1164.all;

LIBRARY work;

ENTITY \32writeenabledflipflop32bit2input\ IS
	PORT
	(
		WriteEnable :  IN  STD_LOGIC;
		ClockInput :  IN  STD_LOGIC;
		Input1 :  IN  STD_LOGIC_VECTOR(31 DOWNTO 0);
		Input2 :  IN  STD_LOGIC_VECTOR(31 DOWNTO 0);
		Selector1 :  IN  STD_LOGIC_VECTOR(0 TO 4);
		Selector2 :  IN  STD_LOGIC_VECTOR(0 TO 4);
		ResultPin1 :  OUT  STD_LOGIC_VECTOR(31 DOWNTO 0);
		ResultPin2 :  OUT  STD_LOGIC_VECTOR(31 DOWNTO 0)
	);
END \32writeenabledflipflop32bit2input\;

ARCHITECTURE bdf_type OF \32writeenabledflipflop32bit2input\ IS

COMPONENT mux32_32bit
	PORT(Input00 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 Input01 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 Input02 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 Input03 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 Input04 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 Input05 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 Input06 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 Input07 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 Input08 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 Input09 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 Input10 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 Input11 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 Input12 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 Input13 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 Input14 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 Input15 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 Input16 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 Input17 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 Input18 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 Input19 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 Input20 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 Input21 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 Input22 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 Input23 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 Input24 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 Input25 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 Input26 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 Input27 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 Input28 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 Input29 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 Input30 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 Input31 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 Selector : IN STD_LOGIC_VECTOR(4 DOWNTO 0);
		 ResultPin : OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
	);
END COMPONENT;

COMPONENT writeenabledflipflop32bit
	PORT(WriteEnable : IN STD_LOGIC;
		 ClockInput : IN STD_LOGIC;
		 Input : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 OutputRes : OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
	);
END COMPONENT;

COMPONENT and5_1bit
	PORT(Input1 : IN STD_LOGIC;
		 Input2 : IN STD_LOGIC;
		 Input3 : IN STD_LOGIC;
		 Input5 : IN STD_LOGIC;
		 Input4 : IN STD_LOGIC;
		 ResultingPin : OUT STD_LOGIC
	);
END COMPONENT;

SIGNAL	SYNTHESIZED_WIRE_0 :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_1 :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_2 :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_3 :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_4 :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_5 :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_6 :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_7 :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_8 :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_9 :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_10 :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_11 :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_12 :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_13 :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_14 :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_15 :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_16 :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_17 :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_18 :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_19 :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_20 :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_21 :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_22 :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_23 :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_24 :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_25 :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_26 :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_27 :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_28 :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_29 :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_30 :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_31 :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_32 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_33 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_34 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_35 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_36 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_37 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_38 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_39 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_40 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_41 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_42 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_43 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_44 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_45 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_46 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_47 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_48 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_49 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_50 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_51 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_52 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_53 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_54 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_55 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_56 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_57 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_58 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_59 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_60 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_61 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_62 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_63 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_64 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_65 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_66 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_67 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_68 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_69 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_70 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_71 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_72 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_73 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_74 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_75 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_76 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_77 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_78 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_79 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_80 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_81 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_82 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_83 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_84 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_85 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_86 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_87 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_88 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_89 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_90 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_91 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_92 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_93 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_94 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_95 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_96 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_97 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_98 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_99 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_100 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_101 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_102 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_103 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_104 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_105 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_106 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_107 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_108 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_109 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_110 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_111 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_112 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_113 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_114 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_115 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_116 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_117 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_118 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_119 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_120 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_121 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_122 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_123 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_124 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_125 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_126 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_127 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_128 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_129 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_130 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_131 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_132 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_133 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_134 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_135 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_136 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_137 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_138 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_139 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_140 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_141 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_142 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_143 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_144 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_145 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_146 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_147 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_148 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_149 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_150 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_151 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_152 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_153 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_154 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_155 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_156 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_157 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_158 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_159 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_160 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_161 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_162 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_163 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_164 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_165 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_166 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_167 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_168 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_169 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_170 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_171 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_172 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_173 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_174 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_175 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_176 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_177 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_178 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_179 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_180 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_181 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_182 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_183 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_184 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_185 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_186 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_187 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_188 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_189 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_190 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_191 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_192 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_193 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_194 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_195 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_196 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_197 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_198 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_199 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_200 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_201 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_202 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_203 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_204 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_205 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_206 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_207 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_384 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_209 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_211 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_213 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_215 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_217 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_219 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_221 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_223 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_225 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_227 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_229 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_231 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_233 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_235 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_237 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_239 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_241 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_243 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_245 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_247 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_249 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_251 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_253 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_255 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_257 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_259 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_261 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_263 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_265 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_267 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_269 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_271 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_272 :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_273 :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_274 :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_275 :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_276 :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_277 :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_278 :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_279 :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_280 :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_281 :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_282 :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_283 :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_284 :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_285 :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_286 :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_287 :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_288 :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_289 :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_290 :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_291 :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_292 :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_293 :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_294 :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_295 :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_296 :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_297 :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_298 :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_299 :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_300 :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_301 :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_302 :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_303 :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_304 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_305 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_306 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_307 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_308 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_309 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_310 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_311 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_312 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_313 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_314 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_315 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_316 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_317 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_318 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_319 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_320 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_321 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_322 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_323 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_324 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_325 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_326 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_327 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_328 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_329 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_330 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_331 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_332 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_333 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_334 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_335 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_336 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_337 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_338 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_339 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_340 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_341 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_342 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_343 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_344 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_345 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_346 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_347 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_348 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_349 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_350 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_351 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_352 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_353 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_354 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_355 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_356 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_357 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_358 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_359 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_360 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_361 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_362 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_363 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_364 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_365 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_366 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_367 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_368 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_369 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_370 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_371 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_372 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_373 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_374 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_375 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_376 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_377 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_378 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_379 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_380 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_381 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_382 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_383 :  STD_LOGIC;


BEGIN
SYNTHESIZED_WIRE_384 <= '0';



b2v_inst : mux32_32bit
PORT MAP(Input00 => SYNTHESIZED_WIRE_0,
		 Input01 => SYNTHESIZED_WIRE_1,
		 Input02 => SYNTHESIZED_WIRE_2,
		 Input03 => SYNTHESIZED_WIRE_3,
		 Input04 => SYNTHESIZED_WIRE_4,
		 Input05 => SYNTHESIZED_WIRE_5,
		 Input06 => SYNTHESIZED_WIRE_6,
		 Input07 => SYNTHESIZED_WIRE_7,
		 Input08 => SYNTHESIZED_WIRE_8,
		 Input09 => SYNTHESIZED_WIRE_9,
		 Input10 => SYNTHESIZED_WIRE_10,
		 Input11 => SYNTHESIZED_WIRE_11,
		 Input12 => SYNTHESIZED_WIRE_12,
		 Input13 => SYNTHESIZED_WIRE_13,
		 Input14 => SYNTHESIZED_WIRE_14,
		 Input15 => SYNTHESIZED_WIRE_15,
		 Input16 => SYNTHESIZED_WIRE_16,
		 Input17 => SYNTHESIZED_WIRE_17,
		 Input18 => SYNTHESIZED_WIRE_18,
		 Input19 => SYNTHESIZED_WIRE_19,
		 Input20 => SYNTHESIZED_WIRE_20,
		 Input21 => SYNTHESIZED_WIRE_21,
		 Input22 => SYNTHESIZED_WIRE_22,
		 Input23 => SYNTHESIZED_WIRE_23,
		 Input24 => SYNTHESIZED_WIRE_24,
		 Input25 => SYNTHESIZED_WIRE_25,
		 Input26 => SYNTHESIZED_WIRE_26,
		 Input27 => SYNTHESIZED_WIRE_27,
		 Input28 => SYNTHESIZED_WIRE_28,
		 Input29 => SYNTHESIZED_WIRE_29,
		 Input30 => SYNTHESIZED_WIRE_30,
		 Input31 => SYNTHESIZED_WIRE_31,
		 Selector => Selector1,
		 ResultPin => ResultPin1);


SYNTHESIZED_WIRE_104 <= NOT(Selector1(4));



SYNTHESIZED_WIRE_100 <= NOT(Selector1(4));



SYNTHESIZED_WIRE_318 <= NOT(Selector2(0));



SYNTHESIZED_WIRE_319 <= NOT(Selector2(4));



SYNTHESIZED_WIRE_320 <= NOT(Selector2(3));



SYNTHESIZED_WIRE_321 <= NOT(Selector2(1));



SYNTHESIZED_WIRE_322 <= NOT(Selector2(4));



SYNTHESIZED_WIRE_323 <= NOT(Selector2(3));



SYNTHESIZED_WIRE_324 <= NOT(Selector2(0));



SYNTHESIZED_WIRE_325 <= NOT(Selector2(4));



SYNTHESIZED_WIRE_326 <= NOT(Selector2(3));



SYNTHESIZED_WIRE_327 <= NOT(Selector2(4));



SYNTHESIZED_WIRE_101 <= NOT(Selector1(3));



SYNTHESIZED_WIRE_328 <= NOT(Selector2(2));



SYNTHESIZED_WIRE_329 <= NOT(Selector2(1));



SYNTHESIZED_WIRE_330 <= NOT(Selector2(0));



SYNTHESIZED_WIRE_64 <= SYNTHESIZED_WIRE_32 AND ClockInput;


SYNTHESIZED_WIRE_65 <= SYNTHESIZED_WIRE_33 AND ClockInput;


SYNTHESIZED_WIRE_66 <= SYNTHESIZED_WIRE_34 AND ClockInput;


SYNTHESIZED_WIRE_67 <= SYNTHESIZED_WIRE_35 AND ClockInput;


SYNTHESIZED_WIRE_68 <= SYNTHESIZED_WIRE_36 AND ClockInput;


SYNTHESIZED_WIRE_69 <= SYNTHESIZED_WIRE_37 AND ClockInput;


SYNTHESIZED_WIRE_70 <= SYNTHESIZED_WIRE_38 AND ClockInput;


SYNTHESIZED_WIRE_102 <= NOT(Selector1(2));



SYNTHESIZED_WIRE_71 <= SYNTHESIZED_WIRE_39 AND ClockInput;


SYNTHESIZED_WIRE_72 <= SYNTHESIZED_WIRE_40 AND ClockInput;


SYNTHESIZED_WIRE_73 <= SYNTHESIZED_WIRE_41 AND ClockInput;


SYNTHESIZED_WIRE_74 <= SYNTHESIZED_WIRE_42 AND ClockInput;


SYNTHESIZED_WIRE_75 <= SYNTHESIZED_WIRE_43 AND ClockInput;


SYNTHESIZED_WIRE_76 <= SYNTHESIZED_WIRE_44 AND ClockInput;


SYNTHESIZED_WIRE_77 <= SYNTHESIZED_WIRE_45 AND ClockInput;


SYNTHESIZED_WIRE_78 <= SYNTHESIZED_WIRE_46 AND ClockInput;


SYNTHESIZED_WIRE_79 <= SYNTHESIZED_WIRE_47 AND ClockInput;


SYNTHESIZED_WIRE_80 <= SYNTHESIZED_WIRE_48 AND ClockInput;


SYNTHESIZED_WIRE_103 <= NOT(Selector1(0));



SYNTHESIZED_WIRE_81 <= SYNTHESIZED_WIRE_49 AND ClockInput;


SYNTHESIZED_WIRE_82 <= SYNTHESIZED_WIRE_50 AND ClockInput;


SYNTHESIZED_WIRE_83 <= SYNTHESIZED_WIRE_51 AND ClockInput;


SYNTHESIZED_WIRE_84 <= SYNTHESIZED_WIRE_52 AND ClockInput;


SYNTHESIZED_WIRE_85 <= SYNTHESIZED_WIRE_53 AND ClockInput;


SYNTHESIZED_WIRE_86 <= SYNTHESIZED_WIRE_54 AND ClockInput;


SYNTHESIZED_WIRE_87 <= SYNTHESIZED_WIRE_55 AND ClockInput;


SYNTHESIZED_WIRE_88 <= SYNTHESIZED_WIRE_56 AND ClockInput;


SYNTHESIZED_WIRE_89 <= SYNTHESIZED_WIRE_57 AND ClockInput;


SYNTHESIZED_WIRE_90 <= SYNTHESIZED_WIRE_58 AND ClockInput;


SYNTHESIZED_WIRE_109 <= NOT(Selector1(4));



SYNTHESIZED_WIRE_91 <= SYNTHESIZED_WIRE_59 AND ClockInput;


SYNTHESIZED_WIRE_92 <= SYNTHESIZED_WIRE_60 AND ClockInput;


SYNTHESIZED_WIRE_93 <= SYNTHESIZED_WIRE_61 AND ClockInput;


SYNTHESIZED_WIRE_94 <= SYNTHESIZED_WIRE_62 AND ClockInput;


SYNTHESIZED_WIRE_95 <= SYNTHESIZED_WIRE_63 AND ClockInput;


b2v_inst145 : writeenabledflipflop32bit
PORT MAP(WriteEnable => WriteEnable,
		 ClockInput => SYNTHESIZED_WIRE_64,
		 Input => Input1,
		 OutputRes => SYNTHESIZED_WIRE_0);


b2v_inst146 : writeenabledflipflop32bit
PORT MAP(WriteEnable => WriteEnable,
		 ClockInput => SYNTHESIZED_WIRE_65,
		 Input => Input1,
		 OutputRes => SYNTHESIZED_WIRE_1);


b2v_inst147 : writeenabledflipflop32bit
PORT MAP(WriteEnable => WriteEnable,
		 ClockInput => SYNTHESIZED_WIRE_66,
		 Input => Input1,
		 OutputRes => SYNTHESIZED_WIRE_2);


b2v_inst148 : writeenabledflipflop32bit
PORT MAP(WriteEnable => WriteEnable,
		 ClockInput => SYNTHESIZED_WIRE_67,
		 Input => Input1,
		 OutputRes => SYNTHESIZED_WIRE_3);


b2v_inst149 : writeenabledflipflop32bit
PORT MAP(WriteEnable => WriteEnable,
		 ClockInput => SYNTHESIZED_WIRE_68,
		 Input => Input1,
		 OutputRes => SYNTHESIZED_WIRE_4);


SYNTHESIZED_WIRE_110 <= NOT(Selector1(3));



b2v_inst150 : writeenabledflipflop32bit
PORT MAP(WriteEnable => WriteEnable,
		 ClockInput => SYNTHESIZED_WIRE_69,
		 Input => Input1,
		 OutputRes => SYNTHESIZED_WIRE_5);


b2v_inst151 : writeenabledflipflop32bit
PORT MAP(WriteEnable => WriteEnable,
		 ClockInput => SYNTHESIZED_WIRE_70,
		 Input => Input1,
		 OutputRes => SYNTHESIZED_WIRE_6);


b2v_inst152 : writeenabledflipflop32bit
PORT MAP(WriteEnable => WriteEnable,
		 ClockInput => SYNTHESIZED_WIRE_71,
		 Input => Input1,
		 OutputRes => SYNTHESIZED_WIRE_7);


b2v_inst153 : writeenabledflipflop32bit
PORT MAP(WriteEnable => WriteEnable,
		 ClockInput => SYNTHESIZED_WIRE_72,
		 Input => Input1,
		 OutputRes => SYNTHESIZED_WIRE_8);


b2v_inst154 : writeenabledflipflop32bit
PORT MAP(WriteEnable => WriteEnable,
		 ClockInput => SYNTHESIZED_WIRE_73,
		 Input => Input1,
		 OutputRes => SYNTHESIZED_WIRE_9);


b2v_inst155 : writeenabledflipflop32bit
PORT MAP(WriteEnable => WriteEnable,
		 ClockInput => SYNTHESIZED_WIRE_74,
		 Input => Input1,
		 OutputRes => SYNTHESIZED_WIRE_10);


b2v_inst156 : writeenabledflipflop32bit
PORT MAP(WriteEnable => WriteEnable,
		 ClockInput => SYNTHESIZED_WIRE_75,
		 Input => Input1,
		 OutputRes => SYNTHESIZED_WIRE_11);


b2v_inst157 : writeenabledflipflop32bit
PORT MAP(WriteEnable => WriteEnable,
		 ClockInput => SYNTHESIZED_WIRE_76,
		 Input => Input1,
		 OutputRes => SYNTHESIZED_WIRE_12);


b2v_inst158 : writeenabledflipflop32bit
PORT MAP(WriteEnable => WriteEnable,
		 ClockInput => SYNTHESIZED_WIRE_77,
		 Input => Input1,
		 OutputRes => SYNTHESIZED_WIRE_13);


b2v_inst159 : writeenabledflipflop32bit
PORT MAP(WriteEnable => WriteEnable,
		 ClockInput => SYNTHESIZED_WIRE_78,
		 Input => Input1,
		 OutputRes => SYNTHESIZED_WIRE_14);


SYNTHESIZED_WIRE_111 <= NOT(Selector1(2));



b2v_inst160 : writeenabledflipflop32bit
PORT MAP(WriteEnable => WriteEnable,
		 ClockInput => SYNTHESIZED_WIRE_79,
		 Input => Input1,
		 OutputRes => SYNTHESIZED_WIRE_15);


b2v_inst161 : writeenabledflipflop32bit
PORT MAP(WriteEnable => WriteEnable,
		 ClockInput => SYNTHESIZED_WIRE_80,
		 Input => Input1,
		 OutputRes => SYNTHESIZED_WIRE_16);


b2v_inst162 : writeenabledflipflop32bit
PORT MAP(WriteEnable => WriteEnable,
		 ClockInput => SYNTHESIZED_WIRE_81,
		 Input => Input1,
		 OutputRes => SYNTHESIZED_WIRE_17);


b2v_inst163 : writeenabledflipflop32bit
PORT MAP(WriteEnable => WriteEnable,
		 ClockInput => SYNTHESIZED_WIRE_82,
		 Input => Input1,
		 OutputRes => SYNTHESIZED_WIRE_18);


b2v_inst164 : writeenabledflipflop32bit
PORT MAP(WriteEnable => WriteEnable,
		 ClockInput => SYNTHESIZED_WIRE_83,
		 Input => Input1,
		 OutputRes => SYNTHESIZED_WIRE_19);


b2v_inst165 : writeenabledflipflop32bit
PORT MAP(WriteEnable => WriteEnable,
		 ClockInput => SYNTHESIZED_WIRE_84,
		 Input => Input1,
		 OutputRes => SYNTHESIZED_WIRE_20);


b2v_inst166 : writeenabledflipflop32bit
PORT MAP(WriteEnable => WriteEnable,
		 ClockInput => SYNTHESIZED_WIRE_85,
		 Input => Input1,
		 OutputRes => SYNTHESIZED_WIRE_21);


b2v_inst167 : writeenabledflipflop32bit
PORT MAP(WriteEnable => WriteEnable,
		 ClockInput => SYNTHESIZED_WIRE_86,
		 Input => Input1,
		 OutputRes => SYNTHESIZED_WIRE_22);


b2v_inst168 : writeenabledflipflop32bit
PORT MAP(WriteEnable => WriteEnable,
		 ClockInput => SYNTHESIZED_WIRE_87,
		 Input => Input1,
		 OutputRes => SYNTHESIZED_WIRE_23);


b2v_inst169 : writeenabledflipflop32bit
PORT MAP(WriteEnable => WriteEnable,
		 ClockInput => SYNTHESIZED_WIRE_88,
		 Input => Input1,
		 OutputRes => SYNTHESIZED_WIRE_24);


SYNTHESIZED_WIRE_117 <= NOT(Selector1(4));



b2v_inst170 : writeenabledflipflop32bit
PORT MAP(WriteEnable => WriteEnable,
		 ClockInput => SYNTHESIZED_WIRE_89,
		 Input => Input1,
		 OutputRes => SYNTHESIZED_WIRE_25);


b2v_inst171 : writeenabledflipflop32bit
PORT MAP(WriteEnable => WriteEnable,
		 ClockInput => SYNTHESIZED_WIRE_90,
		 Input => Input1,
		 OutputRes => SYNTHESIZED_WIRE_26);


b2v_inst172 : writeenabledflipflop32bit
PORT MAP(WriteEnable => WriteEnable,
		 ClockInput => SYNTHESIZED_WIRE_91,
		 Input => Input1,
		 OutputRes => SYNTHESIZED_WIRE_27);


b2v_inst173 : writeenabledflipflop32bit
PORT MAP(WriteEnable => WriteEnable,
		 ClockInput => SYNTHESIZED_WIRE_92,
		 Input => Input1,
		 OutputRes => SYNTHESIZED_WIRE_28);


b2v_inst174 : writeenabledflipflop32bit
PORT MAP(WriteEnable => WriteEnable,
		 ClockInput => SYNTHESIZED_WIRE_93,
		 Input => Input1,
		 OutputRes => SYNTHESIZED_WIRE_29);


b2v_inst175 : writeenabledflipflop32bit
PORT MAP(WriteEnable => WriteEnable,
		 ClockInput => SYNTHESIZED_WIRE_94,
		 Input => Input1,
		 OutputRes => SYNTHESIZED_WIRE_30);


b2v_inst176 : writeenabledflipflop32bit
PORT MAP(WriteEnable => WriteEnable,
		 ClockInput => SYNTHESIZED_WIRE_95,
		 Input => Input1,
		 OutputRes => SYNTHESIZED_WIRE_31);


SYNTHESIZED_WIRE_331 <= NOT(Selector2(4));



SYNTHESIZED_WIRE_332 <= NOT(Selector2(2));



SYNTHESIZED_WIRE_333 <= NOT(Selector2(1));



SYNTHESIZED_WIRE_118 <= NOT(Selector1(3));



SYNTHESIZED_WIRE_376 <= NOT(Selector2(4));



SYNTHESIZED_WIRE_377 <= NOT(Selector2(2));



SYNTHESIZED_WIRE_378 <= NOT(Selector2(0));



b2v_inst183 : and5_1bit
PORT MAP(Input1 => SYNTHESIZED_WIRE_96,
		 Input2 => SYNTHESIZED_WIRE_97,
		 Input3 => SYNTHESIZED_WIRE_98,
		 Input5 => SYNTHESIZED_WIRE_99,
		 Input4 => Selector1(0),
		 ResultingPin => SYNTHESIZED_WIRE_33);


b2v_inst184 : and5_1bit
PORT MAP(Input1 => SYNTHESIZED_WIRE_100,
		 Input2 => SYNTHESIZED_WIRE_101,
		 Input3 => SYNTHESIZED_WIRE_102,
		 Input5 => Selector1(1),
		 Input4 => SYNTHESIZED_WIRE_103,
		 ResultingPin => SYNTHESIZED_WIRE_34);


b2v_inst185 : and5_1bit
PORT MAP(Input1 => SYNTHESIZED_WIRE_104,
		 Input2 => SYNTHESIZED_WIRE_105,
		 Input3 => SYNTHESIZED_WIRE_106,
		 Input5 => SYNTHESIZED_WIRE_107,
		 Input4 => SYNTHESIZED_WIRE_108,
		 ResultingPin => SYNTHESIZED_WIRE_32);


b2v_inst186 : and5_1bit
PORT MAP(Input1 => SYNTHESIZED_WIRE_109,
		 Input2 => SYNTHESIZED_WIRE_110,
		 Input3 => SYNTHESIZED_WIRE_111,
		 Input5 => Selector1(1),
		 Input4 => Selector1(0),
		 ResultingPin => SYNTHESIZED_WIRE_35);


b2v_inst187 : and5_1bit
PORT MAP(Input1 => SYNTHESIZED_WIRE_112,
		 Input2 => SYNTHESIZED_WIRE_113,
		 Input3 => Selector1(2),
		 Input5 => Selector1(1),
		 Input4 => SYNTHESIZED_WIRE_114,
		 ResultingPin => SYNTHESIZED_WIRE_38);


b2v_inst188 : and5_1bit
PORT MAP(Input1 => SYNTHESIZED_WIRE_115,
		 Input2 => SYNTHESIZED_WIRE_116,
		 Input3 => Selector1(2),
		 Input5 => Selector1(1),
		 Input4 => Selector1(0),
		 ResultingPin => SYNTHESIZED_WIRE_39);


b2v_inst189 : and5_1bit
PORT MAP(Input1 => SYNTHESIZED_WIRE_117,
		 Input2 => SYNTHESIZED_WIRE_118,
		 Input3 => Selector1(2),
		 Input5 => SYNTHESIZED_WIRE_119,
		 Input4 => SYNTHESIZED_WIRE_120,
		 ResultingPin => SYNTHESIZED_WIRE_36);


SYNTHESIZED_WIRE_119 <= NOT(Selector1(1));



b2v_inst190 : and5_1bit
PORT MAP(Input1 => SYNTHESIZED_WIRE_121,
		 Input2 => SYNTHESIZED_WIRE_122,
		 Input3 => Selector1(2),
		 Input5 => SYNTHESIZED_WIRE_123,
		 Input4 => Selector1(0),
		 ResultingPin => SYNTHESIZED_WIRE_37);


b2v_inst191 : and5_1bit
PORT MAP(Input1 => SYNTHESIZED_WIRE_124,
		 Input2 => Selector1(3),
		 Input3 => SYNTHESIZED_WIRE_125,
		 Input5 => SYNTHESIZED_WIRE_126,
		 Input4 => SYNTHESIZED_WIRE_127,
		 ResultingPin => SYNTHESIZED_WIRE_40);


b2v_inst192 : and5_1bit
PORT MAP(Input1 => SYNTHESIZED_WIRE_128,
		 Input2 => Selector1(3),
		 Input3 => SYNTHESIZED_WIRE_129,
		 Input5 => SYNTHESIZED_WIRE_130,
		 Input4 => Selector1(0),
		 ResultingPin => SYNTHESIZED_WIRE_41);


b2v_inst193 : and5_1bit
PORT MAP(Input1 => SYNTHESIZED_WIRE_131,
		 Input2 => Selector1(3),
		 Input3 => SYNTHESIZED_WIRE_132,
		 Input5 => Selector1(1),
		 Input4 => SYNTHESIZED_WIRE_133,
		 ResultingPin => SYNTHESIZED_WIRE_42);


b2v_inst194 : and5_1bit
PORT MAP(Input1 => SYNTHESIZED_WIRE_134,
		 Input2 => Selector1(3),
		 Input3 => SYNTHESIZED_WIRE_135,
		 Input5 => Selector1(1),
		 Input4 => Selector1(0),
		 ResultingPin => SYNTHESIZED_WIRE_43);


b2v_inst195 : and5_1bit
PORT MAP(Input1 => SYNTHESIZED_WIRE_136,
		 Input2 => Selector1(3),
		 Input3 => Selector1(2),
		 Input5 => SYNTHESIZED_WIRE_137,
		 Input4 => SYNTHESIZED_WIRE_138,
		 ResultingPin => SYNTHESIZED_WIRE_44);


b2v_inst196 : and5_1bit
PORT MAP(Input1 => SYNTHESIZED_WIRE_139,
		 Input2 => Selector1(3),
		 Input3 => Selector1(2),
		 Input5 => SYNTHESIZED_WIRE_140,
		 Input4 => Selector1(0),
		 ResultingPin => SYNTHESIZED_WIRE_45);


b2v_inst197 : and5_1bit
PORT MAP(Input1 => SYNTHESIZED_WIRE_141,
		 Input2 => Selector1(3),
		 Input3 => Selector1(2),
		 Input5 => Selector1(1),
		 Input4 => SYNTHESIZED_WIRE_142,
		 ResultingPin => SYNTHESIZED_WIRE_46);


b2v_inst198 : and5_1bit
PORT MAP(Input1 => SYNTHESIZED_WIRE_143,
		 Input2 => Selector1(3),
		 Input3 => Selector1(2),
		 Input5 => Selector1(1),
		 Input4 => Selector1(0),
		 ResultingPin => SYNTHESIZED_WIRE_47);


b2v_inst199 : and5_1bit
PORT MAP(Input1 => Selector1(4),
		 Input2 => SYNTHESIZED_WIRE_144,
		 Input3 => SYNTHESIZED_WIRE_145,
		 Input5 => SYNTHESIZED_WIRE_146,
		 Input4 => SYNTHESIZED_WIRE_147,
		 ResultingPin => SYNTHESIZED_WIRE_48);


SYNTHESIZED_WIRE_105 <= NOT(Selector1(3));



SYNTHESIZED_WIRE_120 <= NOT(Selector1(0));



b2v_inst200 : and5_1bit
PORT MAP(Input1 => Selector1(4),
		 Input2 => SYNTHESIZED_WIRE_148,
		 Input3 => SYNTHESIZED_WIRE_149,
		 Input5 => SYNTHESIZED_WIRE_150,
		 Input4 => Selector1(0),
		 ResultingPin => SYNTHESIZED_WIRE_49);


b2v_inst201 : and5_1bit
PORT MAP(Input1 => Selector1(4),
		 Input2 => SYNTHESIZED_WIRE_151,
		 Input3 => SYNTHESIZED_WIRE_152,
		 Input5 => Selector1(1),
		 Input4 => SYNTHESIZED_WIRE_153,
		 ResultingPin => SYNTHESIZED_WIRE_50);


b2v_inst202 : and5_1bit
PORT MAP(Input1 => Selector1(4),
		 Input2 => SYNTHESIZED_WIRE_154,
		 Input3 => SYNTHESIZED_WIRE_155,
		 Input5 => Selector1(1),
		 Input4 => Selector1(0),
		 ResultingPin => SYNTHESIZED_WIRE_51);


b2v_inst203 : and5_1bit
PORT MAP(Input1 => Selector1(4),
		 Input2 => SYNTHESIZED_WIRE_156,
		 Input3 => Selector1(2),
		 Input5 => SYNTHESIZED_WIRE_157,
		 Input4 => SYNTHESIZED_WIRE_158,
		 ResultingPin => SYNTHESIZED_WIRE_52);


b2v_inst204 : and5_1bit
PORT MAP(Input1 => Selector1(4),
		 Input2 => SYNTHESIZED_WIRE_159,
		 Input3 => Selector1(2),
		 Input5 => SYNTHESIZED_WIRE_160,
		 Input4 => Selector1(0),
		 ResultingPin => SYNTHESIZED_WIRE_53);


b2v_inst205 : and5_1bit
PORT MAP(Input1 => Selector1(4),
		 Input2 => SYNTHESIZED_WIRE_161,
		 Input3 => Selector1(2),
		 Input5 => Selector1(1),
		 Input4 => SYNTHESIZED_WIRE_162,
		 ResultingPin => SYNTHESIZED_WIRE_54);


b2v_inst206 : and5_1bit
PORT MAP(Input1 => Selector1(4),
		 Input2 => SYNTHESIZED_WIRE_163,
		 Input3 => Selector1(2),
		 Input5 => Selector1(1),
		 Input4 => Selector1(0),
		 ResultingPin => SYNTHESIZED_WIRE_55);


b2v_inst207 : and5_1bit
PORT MAP(Input1 => Selector1(4),
		 Input2 => Selector1(3),
		 Input3 => SYNTHESIZED_WIRE_164,
		 Input5 => SYNTHESIZED_WIRE_165,
		 Input4 => SYNTHESIZED_WIRE_166,
		 ResultingPin => SYNTHESIZED_WIRE_56);


b2v_inst208 : and5_1bit
PORT MAP(Input1 => Selector1(4),
		 Input2 => Selector1(3),
		 Input3 => SYNTHESIZED_WIRE_167,
		 Input5 => SYNTHESIZED_WIRE_168,
		 Input4 => Selector1(0),
		 ResultingPin => SYNTHESIZED_WIRE_57);


b2v_inst209 : and5_1bit
PORT MAP(Input1 => Selector1(4),
		 Input2 => Selector1(3),
		 Input3 => SYNTHESIZED_WIRE_169,
		 Input5 => Selector1(1),
		 Input4 => SYNTHESIZED_WIRE_170,
		 ResultingPin => SYNTHESIZED_WIRE_58);


SYNTHESIZED_WIRE_121 <= NOT(Selector1(4));



b2v_inst210 : and5_1bit
PORT MAP(Input1 => Selector1(4),
		 Input2 => Selector1(3),
		 Input3 => SYNTHESIZED_WIRE_171,
		 Input5 => Selector1(1),
		 Input4 => Selector1(0),
		 ResultingPin => SYNTHESIZED_WIRE_59);


b2v_inst211 : and5_1bit
PORT MAP(Input1 => Selector1(4),
		 Input2 => Selector1(3),
		 Input3 => Selector1(2),
		 Input5 => SYNTHESIZED_WIRE_172,
		 Input4 => SYNTHESIZED_WIRE_173,
		 ResultingPin => SYNTHESIZED_WIRE_60);


b2v_inst212 : and5_1bit
PORT MAP(Input1 => Selector1(4),
		 Input2 => Selector1(3),
		 Input3 => Selector1(2),
		 Input5 => SYNTHESIZED_WIRE_174,
		 Input4 => Selector1(0),
		 ResultingPin => SYNTHESIZED_WIRE_61);


b2v_inst213 : and5_1bit
PORT MAP(Input1 => Selector1(4),
		 Input2 => Selector1(3),
		 Input3 => Selector1(2),
		 Input5 => Selector1(1),
		 Input4 => SYNTHESIZED_WIRE_175,
		 ResultingPin => SYNTHESIZED_WIRE_62);


b2v_inst214 : and5_1bit
PORT MAP(Input1 => Selector1(4),
		 Input2 => Selector1(3),
		 Input3 => Selector1(2),
		 Input5 => Selector1(1),
		 Input4 => Selector1(0),
		 ResultingPin => SYNTHESIZED_WIRE_63);


SYNTHESIZED_WIRE_334 <= NOT(Selector2(4));



SYNTHESIZED_WIRE_335 <= NOT(Selector2(2));



SYNTHESIZED_WIRE_336 <= NOT(Selector2(4));



SYNTHESIZED_WIRE_337 <= NOT(Selector2(1));



SYNTHESIZED_WIRE_338 <= NOT(Selector2(0));



SYNTHESIZED_WIRE_122 <= NOT(Selector1(3));



SYNTHESIZED_WIRE_339 <= NOT(Selector2(4));



SYNTHESIZED_WIRE_340 <= NOT(Selector2(1));



SYNTHESIZED_WIRE_341 <= NOT(Selector2(4));



SYNTHESIZED_WIRE_342 <= NOT(Selector2(0));



SYNTHESIZED_WIRE_343 <= NOT(Selector2(4));



SYNTHESIZED_WIRE_344 <= NOT(Selector2(3));



SYNTHESIZED_WIRE_345 <= NOT(Selector2(2));



SYNTHESIZED_WIRE_346 <= NOT(Selector2(1));



SYNTHESIZED_WIRE_347 <= NOT(Selector2(0));



SYNTHESIZED_WIRE_348 <= NOT(Selector2(3));



SYNTHESIZED_WIRE_123 <= NOT(Selector1(1));



SYNTHESIZED_WIRE_349 <= NOT(Selector2(2));



SYNTHESIZED_WIRE_350 <= NOT(Selector2(1));



SYNTHESIZED_WIRE_351 <= NOT(Selector2(3));



SYNTHESIZED_WIRE_352 <= NOT(Selector2(2));



SYNTHESIZED_WIRE_353 <= NOT(Selector2(0));



SYNTHESIZED_WIRE_354 <= NOT(Selector2(3));



SYNTHESIZED_WIRE_355 <= NOT(Selector2(2));



SYNTHESIZED_WIRE_356 <= NOT(Selector2(3));



SYNTHESIZED_WIRE_357 <= NOT(Selector2(1));



SYNTHESIZED_WIRE_358 <= NOT(Selector2(0));



SYNTHESIZED_WIRE_112 <= NOT(Selector1(4));



SYNTHESIZED_WIRE_359 <= NOT(Selector2(3));



SYNTHESIZED_WIRE_360 <= NOT(Selector2(1));



SYNTHESIZED_WIRE_361 <= NOT(Selector2(3));



SYNTHESIZED_WIRE_362 <= NOT(Selector2(0));



SYNTHESIZED_WIRE_363 <= NOT(Selector2(3));



SYNTHESIZED_WIRE_364 <= NOT(Selector2(2));



SYNTHESIZED_WIRE_365 <= NOT(Selector2(1));



SYNTHESIZED_WIRE_366 <= NOT(Selector2(0));



SYNTHESIZED_WIRE_374 <= NOT(Selector2(2));



SYNTHESIZED_WIRE_375 <= NOT(Selector2(1));



SYNTHESIZED_WIRE_113 <= NOT(Selector1(3));



SYNTHESIZED_WIRE_367 <= NOT(Selector2(2));



SYNTHESIZED_WIRE_368 <= NOT(Selector2(0));



SYNTHESIZED_WIRE_369 <= NOT(Selector2(2));



SYNTHESIZED_WIRE_370 <= NOT(Selector2(1));



SYNTHESIZED_WIRE_371 <= NOT(Selector2(0));



SYNTHESIZED_WIRE_372 <= NOT(Selector2(1));



SYNTHESIZED_WIRE_373 <= NOT(Selector2(0));



SYNTHESIZED_WIRE_209 <= SYNTHESIZED_WIRE_176 AND ClockInput;


SYNTHESIZED_WIRE_211 <= SYNTHESIZED_WIRE_177 AND ClockInput;


SYNTHESIZED_WIRE_213 <= SYNTHESIZED_WIRE_178 AND ClockInput;


SYNTHESIZED_WIRE_114 <= NOT(Selector1(0));



SYNTHESIZED_WIRE_215 <= SYNTHESIZED_WIRE_179 AND ClockInput;


SYNTHESIZED_WIRE_217 <= SYNTHESIZED_WIRE_180 AND ClockInput;


SYNTHESIZED_WIRE_219 <= SYNTHESIZED_WIRE_181 AND ClockInput;


SYNTHESIZED_WIRE_221 <= SYNTHESIZED_WIRE_182 AND ClockInput;


SYNTHESIZED_WIRE_223 <= SYNTHESIZED_WIRE_183 AND ClockInput;


SYNTHESIZED_WIRE_225 <= SYNTHESIZED_WIRE_184 AND ClockInput;


SYNTHESIZED_WIRE_227 <= SYNTHESIZED_WIRE_185 AND ClockInput;


SYNTHESIZED_WIRE_229 <= SYNTHESIZED_WIRE_186 AND ClockInput;


SYNTHESIZED_WIRE_231 <= SYNTHESIZED_WIRE_187 AND ClockInput;


SYNTHESIZED_WIRE_233 <= SYNTHESIZED_WIRE_188 AND ClockInput;


SYNTHESIZED_WIRE_115 <= NOT(Selector1(4));



SYNTHESIZED_WIRE_235 <= SYNTHESIZED_WIRE_189 AND ClockInput;


SYNTHESIZED_WIRE_237 <= SYNTHESIZED_WIRE_190 AND ClockInput;


SYNTHESIZED_WIRE_239 <= SYNTHESIZED_WIRE_191 AND ClockInput;


SYNTHESIZED_WIRE_241 <= SYNTHESIZED_WIRE_192 AND ClockInput;


SYNTHESIZED_WIRE_243 <= SYNTHESIZED_WIRE_193 AND ClockInput;


SYNTHESIZED_WIRE_245 <= SYNTHESIZED_WIRE_194 AND ClockInput;


SYNTHESIZED_WIRE_247 <= SYNTHESIZED_WIRE_195 AND ClockInput;


SYNTHESIZED_WIRE_249 <= SYNTHESIZED_WIRE_196 AND ClockInput;


SYNTHESIZED_WIRE_251 <= SYNTHESIZED_WIRE_197 AND ClockInput;


SYNTHESIZED_WIRE_253 <= SYNTHESIZED_WIRE_198 AND ClockInput;


SYNTHESIZED_WIRE_116 <= NOT(Selector1(3));



SYNTHESIZED_WIRE_255 <= SYNTHESIZED_WIRE_199 AND ClockInput;


SYNTHESIZED_WIRE_257 <= SYNTHESIZED_WIRE_200 AND ClockInput;


SYNTHESIZED_WIRE_259 <= SYNTHESIZED_WIRE_201 AND ClockInput;


SYNTHESIZED_WIRE_261 <= SYNTHESIZED_WIRE_202 AND ClockInput;


SYNTHESIZED_WIRE_263 <= SYNTHESIZED_WIRE_203 AND ClockInput;


SYNTHESIZED_WIRE_265 <= SYNTHESIZED_WIRE_204 AND ClockInput;


SYNTHESIZED_WIRE_267 <= SYNTHESIZED_WIRE_205 AND ClockInput;


SYNTHESIZED_WIRE_269 <= SYNTHESIZED_WIRE_206 AND ClockInput;


SYNTHESIZED_WIRE_271 <= SYNTHESIZED_WIRE_207 AND ClockInput;


b2v_inst289 : writeenabledflipflop32bit
PORT MAP(WriteEnable => SYNTHESIZED_WIRE_384,
		 ClockInput => SYNTHESIZED_WIRE_209,
		 Input => Input2,
		 OutputRes => SYNTHESIZED_WIRE_272);


SYNTHESIZED_WIRE_124 <= NOT(Selector1(4));



b2v_inst290 : writeenabledflipflop32bit
PORT MAP(WriteEnable => SYNTHESIZED_WIRE_384,
		 ClockInput => SYNTHESIZED_WIRE_211,
		 Input => Input2,
		 OutputRes => SYNTHESIZED_WIRE_273);


b2v_inst291 : writeenabledflipflop32bit
PORT MAP(WriteEnable => SYNTHESIZED_WIRE_384,
		 ClockInput => SYNTHESIZED_WIRE_213,
		 Input => Input2,
		 OutputRes => SYNTHESIZED_WIRE_274);


b2v_inst292 : writeenabledflipflop32bit
PORT MAP(WriteEnable => SYNTHESIZED_WIRE_384,
		 ClockInput => SYNTHESIZED_WIRE_215,
		 Input => Input2,
		 OutputRes => SYNTHESIZED_WIRE_275);


b2v_inst293 : writeenabledflipflop32bit
PORT MAP(WriteEnable => SYNTHESIZED_WIRE_384,
		 ClockInput => SYNTHESIZED_WIRE_217,
		 Input => Input2,
		 OutputRes => SYNTHESIZED_WIRE_276);


b2v_inst294 : writeenabledflipflop32bit
PORT MAP(WriteEnable => SYNTHESIZED_WIRE_384,
		 ClockInput => SYNTHESIZED_WIRE_219,
		 Input => Input2,
		 OutputRes => SYNTHESIZED_WIRE_277);


b2v_inst295 : writeenabledflipflop32bit
PORT MAP(WriteEnable => SYNTHESIZED_WIRE_384,
		 ClockInput => SYNTHESIZED_WIRE_221,
		 Input => Input2,
		 OutputRes => SYNTHESIZED_WIRE_278);


b2v_inst296 : writeenabledflipflop32bit
PORT MAP(WriteEnable => SYNTHESIZED_WIRE_384,
		 ClockInput => SYNTHESIZED_WIRE_223,
		 Input => Input2,
		 OutputRes => SYNTHESIZED_WIRE_279);


b2v_inst297 : writeenabledflipflop32bit
PORT MAP(WriteEnable => SYNTHESIZED_WIRE_384,
		 ClockInput => SYNTHESIZED_WIRE_225,
		 Input => Input2,
		 OutputRes => SYNTHESIZED_WIRE_280);


b2v_inst298 : writeenabledflipflop32bit
PORT MAP(WriteEnable => SYNTHESIZED_WIRE_384,
		 ClockInput => SYNTHESIZED_WIRE_227,
		 Input => Input2,
		 OutputRes => SYNTHESIZED_WIRE_281);


b2v_inst299 : writeenabledflipflop32bit
PORT MAP(WriteEnable => SYNTHESIZED_WIRE_384,
		 ClockInput => SYNTHESIZED_WIRE_229,
		 Input => Input2,
		 OutputRes => SYNTHESIZED_WIRE_282);


SYNTHESIZED_WIRE_106 <= NOT(Selector1(2));



SYNTHESIZED_WIRE_125 <= NOT(Selector1(2));



b2v_inst300 : writeenabledflipflop32bit
PORT MAP(WriteEnable => SYNTHESIZED_WIRE_384,
		 ClockInput => SYNTHESIZED_WIRE_231,
		 Input => Input2,
		 OutputRes => SYNTHESIZED_WIRE_283);


b2v_inst301 : writeenabledflipflop32bit
PORT MAP(WriteEnable => SYNTHESIZED_WIRE_384,
		 ClockInput => SYNTHESIZED_WIRE_233,
		 Input => Input2,
		 OutputRes => SYNTHESIZED_WIRE_284);


b2v_inst302 : writeenabledflipflop32bit
PORT MAP(WriteEnable => SYNTHESIZED_WIRE_384,
		 ClockInput => SYNTHESIZED_WIRE_235,
		 Input => Input2,
		 OutputRes => SYNTHESIZED_WIRE_285);


b2v_inst303 : writeenabledflipflop32bit
PORT MAP(WriteEnable => SYNTHESIZED_WIRE_384,
		 ClockInput => SYNTHESIZED_WIRE_237,
		 Input => Input2,
		 OutputRes => SYNTHESIZED_WIRE_286);


b2v_inst304 : writeenabledflipflop32bit
PORT MAP(WriteEnable => SYNTHESIZED_WIRE_384,
		 ClockInput => SYNTHESIZED_WIRE_239,
		 Input => Input2,
		 OutputRes => SYNTHESIZED_WIRE_287);


b2v_inst305 : writeenabledflipflop32bit
PORT MAP(WriteEnable => SYNTHESIZED_WIRE_384,
		 ClockInput => SYNTHESIZED_WIRE_241,
		 Input => Input2,
		 OutputRes => SYNTHESIZED_WIRE_288);


b2v_inst306 : writeenabledflipflop32bit
PORT MAP(WriteEnable => SYNTHESIZED_WIRE_384,
		 ClockInput => SYNTHESIZED_WIRE_243,
		 Input => Input2,
		 OutputRes => SYNTHESIZED_WIRE_289);


b2v_inst307 : writeenabledflipflop32bit
PORT MAP(WriteEnable => SYNTHESIZED_WIRE_384,
		 ClockInput => SYNTHESIZED_WIRE_245,
		 Input => Input2,
		 OutputRes => SYNTHESIZED_WIRE_290);


b2v_inst308 : writeenabledflipflop32bit
PORT MAP(WriteEnable => SYNTHESIZED_WIRE_384,
		 ClockInput => SYNTHESIZED_WIRE_247,
		 Input => Input2,
		 OutputRes => SYNTHESIZED_WIRE_291);


b2v_inst309 : writeenabledflipflop32bit
PORT MAP(WriteEnable => SYNTHESIZED_WIRE_384,
		 ClockInput => SYNTHESIZED_WIRE_249,
		 Input => Input2,
		 OutputRes => SYNTHESIZED_WIRE_292);


SYNTHESIZED_WIRE_126 <= NOT(Selector1(1));



b2v_inst310 : writeenabledflipflop32bit
PORT MAP(WriteEnable => SYNTHESIZED_WIRE_384,
		 ClockInput => SYNTHESIZED_WIRE_251,
		 Input => Input2,
		 OutputRes => SYNTHESIZED_WIRE_293);


b2v_inst311 : writeenabledflipflop32bit
PORT MAP(WriteEnable => SYNTHESIZED_WIRE_384,
		 ClockInput => SYNTHESIZED_WIRE_253,
		 Input => Input2,
		 OutputRes => SYNTHESIZED_WIRE_294);


b2v_inst312 : writeenabledflipflop32bit
PORT MAP(WriteEnable => SYNTHESIZED_WIRE_384,
		 ClockInput => SYNTHESIZED_WIRE_255,
		 Input => Input2,
		 OutputRes => SYNTHESIZED_WIRE_295);


b2v_inst313 : writeenabledflipflop32bit
PORT MAP(WriteEnable => SYNTHESIZED_WIRE_384,
		 ClockInput => SYNTHESIZED_WIRE_257,
		 Input => Input2,
		 OutputRes => SYNTHESIZED_WIRE_296);


b2v_inst314 : writeenabledflipflop32bit
PORT MAP(WriteEnable => SYNTHESIZED_WIRE_384,
		 ClockInput => SYNTHESIZED_WIRE_259,
		 Input => Input2,
		 OutputRes => SYNTHESIZED_WIRE_297);


b2v_inst315 : writeenabledflipflop32bit
PORT MAP(WriteEnable => SYNTHESIZED_WIRE_384,
		 ClockInput => SYNTHESIZED_WIRE_261,
		 Input => Input2,
		 OutputRes => SYNTHESIZED_WIRE_298);


b2v_inst316 : writeenabledflipflop32bit
PORT MAP(WriteEnable => SYNTHESIZED_WIRE_384,
		 ClockInput => SYNTHESIZED_WIRE_263,
		 Input => Input2,
		 OutputRes => SYNTHESIZED_WIRE_299);


b2v_inst317 : writeenabledflipflop32bit
PORT MAP(WriteEnable => SYNTHESIZED_WIRE_384,
		 ClockInput => SYNTHESIZED_WIRE_265,
		 Input => Input2,
		 OutputRes => SYNTHESIZED_WIRE_300);


b2v_inst318 : writeenabledflipflop32bit
PORT MAP(WriteEnable => SYNTHESIZED_WIRE_384,
		 ClockInput => SYNTHESIZED_WIRE_267,
		 Input => Input2,
		 OutputRes => SYNTHESIZED_WIRE_301);


b2v_inst319 : writeenabledflipflop32bit
PORT MAP(WriteEnable => SYNTHESIZED_WIRE_384,
		 ClockInput => SYNTHESIZED_WIRE_269,
		 Input => Input2,
		 OutputRes => SYNTHESIZED_WIRE_302);


SYNTHESIZED_WIRE_127 <= NOT(Selector1(0));



b2v_inst320 : writeenabledflipflop32bit
PORT MAP(WriteEnable => SYNTHESIZED_WIRE_384,
		 ClockInput => SYNTHESIZED_WIRE_271,
		 Input => Input2,
		 OutputRes => SYNTHESIZED_WIRE_303);


b2v_inst321 : mux32_32bit
PORT MAP(Input00 => SYNTHESIZED_WIRE_272,
		 Input01 => SYNTHESIZED_WIRE_273,
		 Input02 => SYNTHESIZED_WIRE_274,
		 Input03 => SYNTHESIZED_WIRE_275,
		 Input04 => SYNTHESIZED_WIRE_276,
		 Input05 => SYNTHESIZED_WIRE_277,
		 Input06 => SYNTHESIZED_WIRE_278,
		 Input07 => SYNTHESIZED_WIRE_279,
		 Input08 => SYNTHESIZED_WIRE_280,
		 Input09 => SYNTHESIZED_WIRE_281,
		 Input10 => SYNTHESIZED_WIRE_282,
		 Input11 => SYNTHESIZED_WIRE_283,
		 Input12 => SYNTHESIZED_WIRE_284,
		 Input13 => SYNTHESIZED_WIRE_285,
		 Input14 => SYNTHESIZED_WIRE_286,
		 Input15 => SYNTHESIZED_WIRE_287,
		 Input16 => SYNTHESIZED_WIRE_288,
		 Input17 => SYNTHESIZED_WIRE_289,
		 Input18 => SYNTHESIZED_WIRE_290,
		 Input19 => SYNTHESIZED_WIRE_291,
		 Input20 => SYNTHESIZED_WIRE_292,
		 Input21 => SYNTHESIZED_WIRE_293,
		 Input22 => SYNTHESIZED_WIRE_294,
		 Input23 => SYNTHESIZED_WIRE_295,
		 Input24 => SYNTHESIZED_WIRE_296,
		 Input25 => SYNTHESIZED_WIRE_297,
		 Input26 => SYNTHESIZED_WIRE_298,
		 Input27 => SYNTHESIZED_WIRE_299,
		 Input28 => SYNTHESIZED_WIRE_300,
		 Input29 => SYNTHESIZED_WIRE_301,
		 Input30 => SYNTHESIZED_WIRE_302,
		 Input31 => SYNTHESIZED_WIRE_303,
		 Selector => Selector2,
		 ResultPin => ResultPin2);


b2v_inst322 : and5_1bit
PORT MAP(Input1 => SYNTHESIZED_WIRE_304,
		 Input2 => SYNTHESIZED_WIRE_305,
		 Input3 => SYNTHESIZED_WIRE_306,
		 Input5 => SYNTHESIZED_WIRE_307,
		 Input4 => Selector2(0),
		 ResultingPin => SYNTHESIZED_WIRE_177);


b2v_inst323 : and5_1bit
PORT MAP(Input1 => SYNTHESIZED_WIRE_308,
		 Input2 => SYNTHESIZED_WIRE_309,
		 Input3 => SYNTHESIZED_WIRE_310,
		 Input5 => Selector2(1),
		 Input4 => SYNTHESIZED_WIRE_311,
		 ResultingPin => SYNTHESIZED_WIRE_178);


b2v_inst324 : and5_1bit
PORT MAP(Input1 => SYNTHESIZED_WIRE_312,
		 Input2 => SYNTHESIZED_WIRE_313,
		 Input3 => SYNTHESIZED_WIRE_314,
		 Input5 => Selector2(1),
		 Input4 => Selector2(0),
		 ResultingPin => SYNTHESIZED_WIRE_179);


b2v_inst325 : and5_1bit
PORT MAP(Input1 => SYNTHESIZED_WIRE_315,
		 Input2 => SYNTHESIZED_WIRE_316,
		 Input3 => Selector2(2),
		 Input5 => SYNTHESIZED_WIRE_317,
		 Input4 => SYNTHESIZED_WIRE_318,
		 ResultingPin => SYNTHESIZED_WIRE_180);


b2v_inst326 : and5_1bit
PORT MAP(Input1 => SYNTHESIZED_WIRE_319,
		 Input2 => SYNTHESIZED_WIRE_320,
		 Input3 => Selector2(2),
		 Input5 => SYNTHESIZED_WIRE_321,
		 Input4 => Selector2(0),
		 ResultingPin => SYNTHESIZED_WIRE_181);


b2v_inst327 : and5_1bit
PORT MAP(Input1 => SYNTHESIZED_WIRE_322,
		 Input2 => SYNTHESIZED_WIRE_323,
		 Input3 => Selector2(2),
		 Input5 => Selector2(1),
		 Input4 => SYNTHESIZED_WIRE_324,
		 ResultingPin => SYNTHESIZED_WIRE_182);


b2v_inst328 : and5_1bit
PORT MAP(Input1 => SYNTHESIZED_WIRE_325,
		 Input2 => SYNTHESIZED_WIRE_326,
		 Input3 => Selector2(2),
		 Input5 => Selector2(1),
		 Input4 => Selector2(0),
		 ResultingPin => SYNTHESIZED_WIRE_183);


b2v_inst329 : and5_1bit
PORT MAP(Input1 => SYNTHESIZED_WIRE_327,
		 Input2 => Selector2(3),
		 Input3 => SYNTHESIZED_WIRE_328,
		 Input5 => SYNTHESIZED_WIRE_329,
		 Input4 => SYNTHESIZED_WIRE_330,
		 ResultingPin => SYNTHESIZED_WIRE_184);


SYNTHESIZED_WIRE_128 <= NOT(Selector1(4));



b2v_inst330 : and5_1bit
PORT MAP(Input1 => SYNTHESIZED_WIRE_331,
		 Input2 => Selector2(3),
		 Input3 => SYNTHESIZED_WIRE_332,
		 Input5 => SYNTHESIZED_WIRE_333,
		 Input4 => Selector2(0),
		 ResultingPin => SYNTHESIZED_WIRE_185);


b2v_inst331 : and5_1bit
PORT MAP(Input1 => SYNTHESIZED_WIRE_334,
		 Input2 => Selector2(3),
		 Input3 => SYNTHESIZED_WIRE_335,
		 Input5 => Selector2(1),
		 Input4 => Selector2(0),
		 ResultingPin => SYNTHESIZED_WIRE_187);


b2v_inst332 : and5_1bit
PORT MAP(Input1 => SYNTHESIZED_WIRE_336,
		 Input2 => Selector2(3),
		 Input3 => Selector2(2),
		 Input5 => SYNTHESIZED_WIRE_337,
		 Input4 => SYNTHESIZED_WIRE_338,
		 ResultingPin => SYNTHESIZED_WIRE_188);


b2v_inst333 : and5_1bit
PORT MAP(Input1 => SYNTHESIZED_WIRE_339,
		 Input2 => Selector2(3),
		 Input3 => Selector2(2),
		 Input5 => SYNTHESIZED_WIRE_340,
		 Input4 => Selector2(0),
		 ResultingPin => SYNTHESIZED_WIRE_189);


b2v_inst334 : and5_1bit
PORT MAP(Input1 => SYNTHESIZED_WIRE_341,
		 Input2 => Selector2(3),
		 Input3 => Selector2(2),
		 Input5 => Selector2(1),
		 Input4 => SYNTHESIZED_WIRE_342,
		 ResultingPin => SYNTHESIZED_WIRE_190);


b2v_inst335 : and5_1bit
PORT MAP(Input1 => SYNTHESIZED_WIRE_343,
		 Input2 => Selector2(3),
		 Input3 => Selector2(2),
		 Input5 => Selector2(1),
		 Input4 => Selector2(0),
		 ResultingPin => SYNTHESIZED_WIRE_191);


b2v_inst336 : and5_1bit
PORT MAP(Input1 => Selector2(4),
		 Input2 => SYNTHESIZED_WIRE_344,
		 Input3 => SYNTHESIZED_WIRE_345,
		 Input5 => SYNTHESIZED_WIRE_346,
		 Input4 => SYNTHESIZED_WIRE_347,
		 ResultingPin => SYNTHESIZED_WIRE_192);


b2v_inst337 : and5_1bit
PORT MAP(Input1 => Selector2(4),
		 Input2 => SYNTHESIZED_WIRE_348,
		 Input3 => SYNTHESIZED_WIRE_349,
		 Input5 => SYNTHESIZED_WIRE_350,
		 Input4 => Selector2(0),
		 ResultingPin => SYNTHESIZED_WIRE_193);


b2v_inst338 : and5_1bit
PORT MAP(Input1 => Selector2(4),
		 Input2 => SYNTHESIZED_WIRE_351,
		 Input3 => SYNTHESIZED_WIRE_352,
		 Input5 => Selector2(1),
		 Input4 => SYNTHESIZED_WIRE_353,
		 ResultingPin => SYNTHESIZED_WIRE_194);


b2v_inst339 : and5_1bit
PORT MAP(Input1 => Selector2(4),
		 Input2 => SYNTHESIZED_WIRE_354,
		 Input3 => SYNTHESIZED_WIRE_355,
		 Input5 => Selector2(1),
		 Input4 => Selector2(0),
		 ResultingPin => SYNTHESIZED_WIRE_195);


SYNTHESIZED_WIRE_129 <= NOT(Selector1(2));



b2v_inst340 : and5_1bit
PORT MAP(Input1 => Selector2(4),
		 Input2 => SYNTHESIZED_WIRE_356,
		 Input3 => Selector2(2),
		 Input5 => SYNTHESIZED_WIRE_357,
		 Input4 => SYNTHESIZED_WIRE_358,
		 ResultingPin => SYNTHESIZED_WIRE_196);


b2v_inst341 : and5_1bit
PORT MAP(Input1 => Selector2(4),
		 Input2 => SYNTHESIZED_WIRE_359,
		 Input3 => Selector2(2),
		 Input5 => SYNTHESIZED_WIRE_360,
		 Input4 => Selector2(0),
		 ResultingPin => SYNTHESIZED_WIRE_197);


b2v_inst342 : and5_1bit
PORT MAP(Input1 => Selector2(4),
		 Input2 => SYNTHESIZED_WIRE_361,
		 Input3 => Selector2(2),
		 Input5 => Selector2(1),
		 Input4 => SYNTHESIZED_WIRE_362,
		 ResultingPin => SYNTHESIZED_WIRE_198);


b2v_inst343 : and5_1bit
PORT MAP(Input1 => Selector2(4),
		 Input2 => SYNTHESIZED_WIRE_363,
		 Input3 => Selector2(2),
		 Input5 => Selector2(1),
		 Input4 => Selector2(0),
		 ResultingPin => SYNTHESIZED_WIRE_199);


b2v_inst344 : and5_1bit
PORT MAP(Input1 => Selector2(4),
		 Input2 => Selector2(3),
		 Input3 => SYNTHESIZED_WIRE_364,
		 Input5 => SYNTHESIZED_WIRE_365,
		 Input4 => SYNTHESIZED_WIRE_366,
		 ResultingPin => SYNTHESIZED_WIRE_200);


b2v_inst345 : and5_1bit
PORT MAP(Input1 => Selector2(4),
		 Input2 => Selector2(3),
		 Input3 => SYNTHESIZED_WIRE_367,
		 Input5 => Selector2(1),
		 Input4 => SYNTHESIZED_WIRE_368,
		 ResultingPin => SYNTHESIZED_WIRE_202);


b2v_inst346 : and5_1bit
PORT MAP(Input1 => Selector2(4),
		 Input2 => Selector2(3),
		 Input3 => SYNTHESIZED_WIRE_369,
		 Input5 => Selector2(1),
		 Input4 => Selector2(0),
		 ResultingPin => SYNTHESIZED_WIRE_203);


b2v_inst347 : and5_1bit
PORT MAP(Input1 => Selector2(4),
		 Input2 => Selector2(3),
		 Input3 => Selector2(2),
		 Input5 => SYNTHESIZED_WIRE_370,
		 Input4 => SYNTHESIZED_WIRE_371,
		 ResultingPin => SYNTHESIZED_WIRE_204);


b2v_inst348 : and5_1bit
PORT MAP(Input1 => Selector2(4),
		 Input2 => Selector2(3),
		 Input3 => Selector2(2),
		 Input5 => SYNTHESIZED_WIRE_372,
		 Input4 => Selector2(0),
		 ResultingPin => SYNTHESIZED_WIRE_205);


b2v_inst349 : and5_1bit
PORT MAP(Input1 => Selector2(4),
		 Input2 => Selector2(3),
		 Input3 => Selector2(2),
		 Input5 => Selector2(1),
		 Input4 => SYNTHESIZED_WIRE_373,
		 ResultingPin => SYNTHESIZED_WIRE_206);


SYNTHESIZED_WIRE_130 <= NOT(Selector1(1));



b2v_inst350 : and5_1bit
PORT MAP(Input1 => Selector2(4),
		 Input2 => Selector2(3),
		 Input3 => Selector2(2),
		 Input5 => Selector2(1),
		 Input4 => Selector2(0),
		 ResultingPin => SYNTHESIZED_WIRE_207);


b2v_inst351 : and5_1bit
PORT MAP(Input1 => Selector2(4),
		 Input2 => Selector2(3),
		 Input3 => SYNTHESIZED_WIRE_374,
		 Input5 => SYNTHESIZED_WIRE_375,
		 Input4 => Selector2(0),
		 ResultingPin => SYNTHESIZED_WIRE_201);


b2v_inst352 : and5_1bit
PORT MAP(Input1 => SYNTHESIZED_WIRE_376,
		 Input2 => Selector2(3),
		 Input3 => SYNTHESIZED_WIRE_377,
		 Input5 => Selector2(1),
		 Input4 => SYNTHESIZED_WIRE_378,
		 ResultingPin => SYNTHESIZED_WIRE_186);


b2v_inst353 : and5_1bit
PORT MAP(Input1 => SYNTHESIZED_WIRE_379,
		 Input2 => SYNTHESIZED_WIRE_380,
		 Input3 => SYNTHESIZED_WIRE_381,
		 Input5 => SYNTHESIZED_WIRE_382,
		 Input4 => SYNTHESIZED_WIRE_383,
		 ResultingPin => SYNTHESIZED_WIRE_176);



SYNTHESIZED_WIRE_131 <= NOT(Selector1(4));



SYNTHESIZED_WIRE_132 <= NOT(Selector1(2));



SYNTHESIZED_WIRE_133 <= NOT(Selector1(0));



SYNTHESIZED_WIRE_134 <= NOT(Selector1(4));



SYNTHESIZED_WIRE_107 <= NOT(Selector1(1));



SYNTHESIZED_WIRE_135 <= NOT(Selector1(2));



SYNTHESIZED_WIRE_136 <= NOT(Selector1(4));



SYNTHESIZED_WIRE_137 <= NOT(Selector1(1));



SYNTHESIZED_WIRE_138 <= NOT(Selector1(0));



SYNTHESIZED_WIRE_139 <= NOT(Selector1(4));



SYNTHESIZED_WIRE_140 <= NOT(Selector1(1));



SYNTHESIZED_WIRE_141 <= NOT(Selector1(4));



SYNTHESIZED_WIRE_142 <= NOT(Selector1(0));



SYNTHESIZED_WIRE_143 <= NOT(Selector1(4));



SYNTHESIZED_WIRE_144 <= NOT(Selector1(3));



SYNTHESIZED_WIRE_108 <= NOT(Selector1(0));



SYNTHESIZED_WIRE_145 <= NOT(Selector1(2));



SYNTHESIZED_WIRE_146 <= NOT(Selector1(1));



SYNTHESIZED_WIRE_147 <= NOT(Selector1(0));



SYNTHESIZED_WIRE_148 <= NOT(Selector1(3));



SYNTHESIZED_WIRE_149 <= NOT(Selector1(2));



SYNTHESIZED_WIRE_150 <= NOT(Selector1(1));



SYNTHESIZED_WIRE_151 <= NOT(Selector1(3));



SYNTHESIZED_WIRE_152 <= NOT(Selector1(2));



SYNTHESIZED_WIRE_153 <= NOT(Selector1(0));



SYNTHESIZED_WIRE_154 <= NOT(Selector1(3));



SYNTHESIZED_WIRE_96 <= NOT(Selector1(4));



SYNTHESIZED_WIRE_155 <= NOT(Selector1(2));



SYNTHESIZED_WIRE_156 <= NOT(Selector1(3));



SYNTHESIZED_WIRE_157 <= NOT(Selector1(1));



SYNTHESIZED_WIRE_158 <= NOT(Selector1(0));



SYNTHESIZED_WIRE_159 <= NOT(Selector1(3));



SYNTHESIZED_WIRE_160 <= NOT(Selector1(1));



SYNTHESIZED_WIRE_161 <= NOT(Selector1(3));



SYNTHESIZED_WIRE_162 <= NOT(Selector1(0));



SYNTHESIZED_WIRE_163 <= NOT(Selector1(3));



SYNTHESIZED_WIRE_164 <= NOT(Selector1(2));



SYNTHESIZED_WIRE_97 <= NOT(Selector1(3));



SYNTHESIZED_WIRE_165 <= NOT(Selector1(1));



SYNTHESIZED_WIRE_166 <= NOT(Selector1(0));



SYNTHESIZED_WIRE_167 <= NOT(Selector1(2));



SYNTHESIZED_WIRE_168 <= NOT(Selector1(1));



SYNTHESIZED_WIRE_169 <= NOT(Selector1(2));



SYNTHESIZED_WIRE_170 <= NOT(Selector1(0));



SYNTHESIZED_WIRE_171 <= NOT(Selector1(2));



SYNTHESIZED_WIRE_172 <= NOT(Selector1(1));



SYNTHESIZED_WIRE_173 <= NOT(Selector1(0));



SYNTHESIZED_WIRE_174 <= NOT(Selector1(1));



SYNTHESIZED_WIRE_98 <= NOT(Selector1(2));



SYNTHESIZED_WIRE_175 <= NOT(Selector1(0));



SYNTHESIZED_WIRE_379 <= NOT(Selector2(4));



SYNTHESIZED_WIRE_380 <= NOT(Selector2(3));



SYNTHESIZED_WIRE_381 <= NOT(Selector2(2));



SYNTHESIZED_WIRE_382 <= NOT(Selector2(1));



SYNTHESIZED_WIRE_383 <= NOT(Selector2(0));



SYNTHESIZED_WIRE_304 <= NOT(Selector2(4));



SYNTHESIZED_WIRE_305 <= NOT(Selector2(3));



SYNTHESIZED_WIRE_306 <= NOT(Selector2(2));



SYNTHESIZED_WIRE_307 <= NOT(Selector2(1));



SYNTHESIZED_WIRE_99 <= NOT(Selector1(1));



SYNTHESIZED_WIRE_308 <= NOT(Selector2(4));



SYNTHESIZED_WIRE_309 <= NOT(Selector2(3));



SYNTHESIZED_WIRE_310 <= NOT(Selector2(2));



SYNTHESIZED_WIRE_311 <= NOT(Selector2(0));



SYNTHESIZED_WIRE_312 <= NOT(Selector2(4));



SYNTHESIZED_WIRE_313 <= NOT(Selector2(3));



SYNTHESIZED_WIRE_314 <= NOT(Selector2(2));



SYNTHESIZED_WIRE_315 <= NOT(Selector2(4));



SYNTHESIZED_WIRE_316 <= NOT(Selector2(3));



SYNTHESIZED_WIRE_317 <= NOT(Selector2(1));



END bdf_type;